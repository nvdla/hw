// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_NVDLA_SDP_CORE_Y_idx.v

module SDP_Y_IDX_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_IDX_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module SDP_Y_IDX_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_IDX_mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module SDP_Y_IDX_mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> ../td_ccore_solutions/leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-183
//  Generated date: Tue Mar  7 18:15:16 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_IDX_leading_sign_32_0
// ------------------------------------------------------------------


module SDP_Y_IDX_leading_sign_32_0 (
  mantissa, rtn
);
  input [31:0] mantissa;
  output [5:0] rtn;


  // Interconnect Declarations
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1;
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;

  wire[4:0] IntLeadZero_32U_leading_sign_32_0_rtn_IntLeadZero_32U_leading_sign_32_0_rtn_and_nl;
  wire[0:0] IntLeadZero_32U_leading_sign_32_0_rtn_and_119_nl;
  wire[0:0] IntLeadZero_32U_leading_sign_32_0_rtn_and_117_nl;
  wire[0:0] IntLeadZero_32U_leading_sign_32_0_rtn_and_124_nl;
  wire[0:0] IntLeadZero_32U_leading_sign_32_0_rtn_and_127_nl;
  wire[0:0] IntLeadZero_32U_leading_sign_32_0_rtn_not_nl;

  // Interconnect Declarations for Component Instantiations 
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[29:28]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[31:30]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[27:26]!=2'b00));
  assign c_h_1_2 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[25:24]==2'b00)
      & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[21:20]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[23:22]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[19:18]!=2'b00));
  assign c_h_1_5 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[17:16]==2'b00)
      & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[13:12]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[15:14]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1 = ~((mantissa[11:10]!=2'b00));
  assign c_h_1_9 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3 = (mantissa[9:8]==2'b00)
      & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2 = ~((mantissa[5:4]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1 = ~((mantissa[7:6]!=2'b00));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1 = ~((mantissa[3:2]!=2'b00));
  assign c_h_1_12 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5 = (mantissa[1:0]==2'b00)
      & IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1 & c_h_1_12 & c_h_1_13
      & c_h_1_14;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_119_nl = c_h_1_6 & (c_h_1_13 |
      (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_117_nl = c_h_1_2 & (c_h_1_5 |
      (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3)) & (~((~(c_h_1_9
      & (c_h_1_12 | (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_124_nl = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1
      | (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2)) & (~((~(IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1
      & (IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1 | (~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_127_nl = (~((mantissa[31]) | (~((mantissa[30:29]!=2'b01)))))
      & (~(((mantissa[27]) | (~((mantissa[26:25]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[23])
      | (~((mantissa[22:21]!=2'b01))))) & (~(((mantissa[19]) | (~((mantissa[18:17]!=2'b01))))
      & c_h_1_5)))) & c_h_1_6)) & (~((~((~((mantissa[15]) | (~((mantissa[14:13]!=2'b01)))))
      & (~(((mantissa[11]) | (~((mantissa[10:9]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[7])
      | (~((mantissa[6:5]!=2'b01))))) & (~(((mantissa[3]) | (~((mantissa[2:1]!=2'b01))))
      & c_h_1_12)))) & c_h_1_13)))) & c_h_1_14));
  assign IntLeadZero_32U_leading_sign_32_0_rtn_not_nl = ~ IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_IntLeadZero_32U_leading_sign_32_0_rtn_and_nl
      = MUX_v_5_2_2(5'b00000, ({c_h_1_14 , (IntLeadZero_32U_leading_sign_32_0_rtn_and_119_nl)
      , (IntLeadZero_32U_leading_sign_32_0_rtn_and_117_nl) , (IntLeadZero_32U_leading_sign_32_0_rtn_and_124_nl)
      , (IntLeadZero_32U_leading_sign_32_0_rtn_and_127_nl)}), (IntLeadZero_32U_leading_sign_32_0_rtn_not_nl));
  assign rtn = {IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5 , (IntLeadZero_32U_leading_sign_32_0_rtn_IntLeadZero_32U_leading_sign_32_0_rtn_and_nl)};

  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction

endmodule




//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v4.v 
module SDP_Y_IDX_mgc_shift_bl_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SIGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v 
module SDP_Y_IDX_mgc_shift_l_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v4.v 
module SDP_Y_IDX_mgc_shift_br_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> ../td_ccore_solutions/leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-136
//  Generated date: Fri Jun 16 21:48:25 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_IDX_leading_sign_49_0
// ------------------------------------------------------------------


module SDP_Y_IDX_leading_sign_49_0 (
  mantissa, rtn
);
  input [48:0] mantissa;
  output [5:0] rtn;


  // Interconnect Declarations
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_22;
  wire c_h_1_23;

  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[42:41]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[34:33]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = (mantissa[26:25]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = (mantissa[18:17]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 & c_h_1_12 & c_h_1_13;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = (mantissa[10:9]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = (mantissa[2:1]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (c_h_1_22
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = c_h_1_6 & (c_h_1_13 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4)) & (~((~(c_h_1_21
      & (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4))) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = c_h_1_2 & (c_h_1_5 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3)) & (~((~(c_h_1_9
      & (c_h_1_12 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~(((~(c_h_1_17 & (c_h_1_20 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2)) & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~(((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2)))) & c_h_1_21))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl
      = ((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01))))) & (~(((mantissa[44])
      | (~((mantissa[43:42]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))))
      & (~(((mantissa[36]) | (~((mantissa[35:34]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01))))) & (~(((mantissa[28])
      | (~((mantissa[27:26]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))))
      & (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~(((~((~((mantissa[16]) | (~((mantissa[15:14]!=2'b01))))) &
      (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[8])
      | (~((mantissa[7:6]!=2'b01))))) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)))) | c_h_1_22) & c_h_1_23))) | ((~ (mantissa[0]))
      & c_h_1_22 & c_h_1_23);
  assign rtn = {c_h_1_23 , (IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl)};
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-207
//  Generated date: Tue Jul  4 14:16:37 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_IDX_chn_lut_out_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_IDX_chn_lut_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_IDX_chn_lut_in_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_IDX_chn_lut_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_staller
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_lut_in_rsci_wen_comp, core_wten,
      chn_lut_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_lut_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_lut_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_lut_in_rsci_wen_comp & chn_lut_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_dp
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_out_rsci_oswt, chn_lut_out_rsci_bawt,
      chn_lut_out_rsci_wen_comp, chn_lut_out_rsci_biwt, chn_lut_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_lut_out_rsci_oswt;
  output chn_lut_out_rsci_bawt;
  output chn_lut_out_rsci_wen_comp;
  input chn_lut_out_rsci_biwt;
  input chn_lut_out_rsci_bdwt;


  // Interconnect Declarations
  reg chn_lut_out_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_lut_out_rsci_bawt = chn_lut_out_rsci_biwt | chn_lut_out_rsci_bcwt;
  assign chn_lut_out_rsci_wen_comp = (~ chn_lut_out_rsci_oswt) | chn_lut_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_lut_out_rsci_bcwt <= ~((~(chn_lut_out_rsci_bcwt | chn_lut_out_rsci_biwt))
          | chn_lut_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_ctrl
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_out_rsci_oswt, core_wen, core_wten, chn_lut_out_rsci_iswt0,
      chn_lut_out_rsci_ld_core_psct, chn_lut_out_rsci_biwt, chn_lut_out_rsci_bdwt,
      chn_lut_out_rsci_ld_core_sct, chn_lut_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_lut_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_lut_out_rsci_iswt0;
  input chn_lut_out_rsci_ld_core_psct;
  output chn_lut_out_rsci_biwt;
  output chn_lut_out_rsci_bdwt;
  output chn_lut_out_rsci_ld_core_sct;
  input chn_lut_out_rsci_vd;


  // Interconnect Declarations
  wire chn_lut_out_rsci_ogwt;
  wire chn_lut_out_rsci_pdswt0;
  reg chn_lut_out_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_lut_out_rsci_pdswt0 = (~ core_wten) & chn_lut_out_rsci_iswt0;
  assign chn_lut_out_rsci_biwt = chn_lut_out_rsci_ogwt & chn_lut_out_rsci_vd;
  assign chn_lut_out_rsci_ogwt = chn_lut_out_rsci_pdswt0 | chn_lut_out_rsci_icwt;
  assign chn_lut_out_rsci_bdwt = chn_lut_out_rsci_oswt & core_wen;
  assign chn_lut_out_rsci_ld_core_sct = chn_lut_out_rsci_ld_core_psct & chn_lut_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_lut_out_rsci_icwt <= ~((~(chn_lut_out_rsci_icwt | chn_lut_out_rsci_pdswt0))
          | chn_lut_out_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_dp
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_in_rsci_oswt, chn_lut_in_rsci_bawt, chn_lut_in_rsci_wen_comp,
      chn_lut_in_rsci_d_mxwt, chn_lut_in_rsci_biwt, chn_lut_in_rsci_bdwt, chn_lut_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_lut_in_rsci_oswt;
  output chn_lut_in_rsci_bawt;
  output chn_lut_in_rsci_wen_comp;
  output [127:0] chn_lut_in_rsci_d_mxwt;
  input chn_lut_in_rsci_biwt;
  input chn_lut_in_rsci_bdwt;
  input [127:0] chn_lut_in_rsci_d;


  // Interconnect Declarations
  reg chn_lut_in_rsci_bcwt;
  reg [127:0] chn_lut_in_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_lut_in_rsci_bawt = chn_lut_in_rsci_biwt | chn_lut_in_rsci_bcwt;
  assign chn_lut_in_rsci_wen_comp = (~ chn_lut_in_rsci_oswt) | chn_lut_in_rsci_bawt;
  assign chn_lut_in_rsci_d_mxwt = MUX_v_128_2_2(chn_lut_in_rsci_d, chn_lut_in_rsci_d_bfwt,
      chn_lut_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_in_rsci_bcwt <= 1'b0;
      chn_lut_in_rsci_d_bfwt <= 128'b0;
    end
    else begin
      chn_lut_in_rsci_bcwt <= ~((~(chn_lut_in_rsci_bcwt | chn_lut_in_rsci_biwt))
          | chn_lut_in_rsci_bdwt);
      chn_lut_in_rsci_d_bfwt <= chn_lut_in_rsci_d_mxwt;
    end
  end

  function [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_ctrl
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_in_rsci_oswt, core_wen, chn_lut_in_rsci_iswt0,
      chn_lut_in_rsci_ld_core_psct, core_wten, chn_lut_in_rsci_biwt, chn_lut_in_rsci_bdwt,
      chn_lut_in_rsci_ld_core_sct, chn_lut_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_lut_in_rsci_oswt;
  input core_wen;
  input chn_lut_in_rsci_iswt0;
  input chn_lut_in_rsci_ld_core_psct;
  input core_wten;
  output chn_lut_in_rsci_biwt;
  output chn_lut_in_rsci_bdwt;
  output chn_lut_in_rsci_ld_core_sct;
  input chn_lut_in_rsci_vd;


  // Interconnect Declarations
  wire chn_lut_in_rsci_ogwt;
  wire chn_lut_in_rsci_pdswt0;
  reg chn_lut_in_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_lut_in_rsci_pdswt0 = (~ core_wten) & chn_lut_in_rsci_iswt0;
  assign chn_lut_in_rsci_biwt = chn_lut_in_rsci_ogwt & chn_lut_in_rsci_vd;
  assign chn_lut_in_rsci_ogwt = chn_lut_in_rsci_pdswt0 | chn_lut_in_rsci_icwt;
  assign chn_lut_in_rsci_bdwt = chn_lut_in_rsci_oswt & core_wen;
  assign chn_lut_in_rsci_ld_core_sct = chn_lut_in_rsci_ld_core_psct & chn_lut_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_lut_in_rsci_icwt <= ~((~(chn_lut_in_rsci_icwt | chn_lut_in_rsci_pdswt0))
          | chn_lut_in_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_out_rsc_z, chn_lut_out_rsc_vz, chn_lut_out_rsc_lz,
      chn_lut_out_rsci_oswt, core_wen, core_wten, chn_lut_out_rsci_iswt0, chn_lut_out_rsci_bawt,
      chn_lut_out_rsci_wen_comp, chn_lut_out_rsci_ld_core_psct, chn_lut_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [323:0] chn_lut_out_rsc_z;
  input chn_lut_out_rsc_vz;
  output chn_lut_out_rsc_lz;
  input chn_lut_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_lut_out_rsci_iswt0;
  output chn_lut_out_rsci_bawt;
  output chn_lut_out_rsci_wen_comp;
  input chn_lut_out_rsci_ld_core_psct;
  input [323:0] chn_lut_out_rsci_d;


  // Interconnect Declarations
  wire chn_lut_out_rsci_biwt;
  wire chn_lut_out_rsci_bdwt;
  wire chn_lut_out_rsci_ld_core_sct;
  wire chn_lut_out_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_IDX_mgc_out_stdreg_wait_v1 #(.rscid(32'sd12),
  .width(32'sd324)) chn_lut_out_rsci (
      .ld(chn_lut_out_rsci_ld_core_sct),
      .vd(chn_lut_out_rsci_vd),
      .d(chn_lut_out_rsci_d),
      .lz(chn_lut_out_rsc_lz),
      .vz(chn_lut_out_rsc_vz),
      .z(chn_lut_out_rsc_z)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_ctrl NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_out_rsci_oswt(chn_lut_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_lut_out_rsci_iswt0(chn_lut_out_rsci_iswt0),
      .chn_lut_out_rsci_ld_core_psct(chn_lut_out_rsci_ld_core_psct),
      .chn_lut_out_rsci_biwt(chn_lut_out_rsci_biwt),
      .chn_lut_out_rsci_bdwt(chn_lut_out_rsci_bdwt),
      .chn_lut_out_rsci_ld_core_sct(chn_lut_out_rsci_ld_core_sct),
      .chn_lut_out_rsci_vd(chn_lut_out_rsci_vd)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_dp NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_chn_lut_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_out_rsci_oswt(chn_lut_out_rsci_oswt),
      .chn_lut_out_rsci_bawt(chn_lut_out_rsci_bawt),
      .chn_lut_out_rsci_wen_comp(chn_lut_out_rsci_wen_comp),
      .chn_lut_out_rsci_biwt(chn_lut_out_rsci_biwt),
      .chn_lut_out_rsci_bdwt(chn_lut_out_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_in_rsc_z, chn_lut_in_rsc_vz, chn_lut_in_rsc_lz,
      chn_lut_in_rsci_oswt, core_wen, chn_lut_in_rsci_iswt0, chn_lut_in_rsci_bawt,
      chn_lut_in_rsci_wen_comp, chn_lut_in_rsci_ld_core_psct, chn_lut_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_lut_in_rsc_z;
  input chn_lut_in_rsc_vz;
  output chn_lut_in_rsc_lz;
  input chn_lut_in_rsci_oswt;
  input core_wen;
  input chn_lut_in_rsci_iswt0;
  output chn_lut_in_rsci_bawt;
  output chn_lut_in_rsci_wen_comp;
  input chn_lut_in_rsci_ld_core_psct;
  output [127:0] chn_lut_in_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_lut_in_rsci_biwt;
  wire chn_lut_in_rsci_bdwt;
  wire chn_lut_in_rsci_ld_core_sct;
  wire chn_lut_in_rsci_vd;
  wire [127:0] chn_lut_in_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_IDX_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd128)) chn_lut_in_rsci (
      .ld(chn_lut_in_rsci_ld_core_sct),
      .vd(chn_lut_in_rsci_vd),
      .d(chn_lut_in_rsci_d),
      .lz(chn_lut_in_rsc_lz),
      .vz(chn_lut_in_rsc_vz),
      .z(chn_lut_in_rsc_z)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_ctrl NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_in_rsci_oswt(chn_lut_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_lut_in_rsci_iswt0(chn_lut_in_rsci_iswt0),
      .chn_lut_in_rsci_ld_core_psct(chn_lut_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_lut_in_rsci_biwt(chn_lut_in_rsci_biwt),
      .chn_lut_in_rsci_bdwt(chn_lut_in_rsci_bdwt),
      .chn_lut_in_rsci_ld_core_sct(chn_lut_in_rsci_ld_core_sct),
      .chn_lut_in_rsci_vd(chn_lut_in_rsci_vd)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_dp NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_chn_lut_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_in_rsci_oswt(chn_lut_in_rsci_oswt),
      .chn_lut_in_rsci_bawt(chn_lut_in_rsci_bawt),
      .chn_lut_in_rsci_wen_comp(chn_lut_in_rsci_wen_comp),
      .chn_lut_in_rsci_d_mxwt(chn_lut_in_rsci_d_mxwt),
      .chn_lut_in_rsci_biwt(chn_lut_in_rsci_biwt),
      .chn_lut_in_rsci_bdwt(chn_lut_in_rsci_bdwt),
      .chn_lut_in_rsci_d(chn_lut_in_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx_core
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx_core (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_in_rsc_z, chn_lut_in_rsc_vz, chn_lut_in_rsc_lz,
      cfg_lut_le_start_rsc_z, cfg_lut_lo_start_rsc_z, cfg_lut_le_index_offset_rsc_z,
      cfg_lut_le_index_select_rsc_z, cfg_lut_lo_index_select_rsc_z, cfg_lut_le_function_rsc_z,
      cfg_lut_uflow_priority_rsc_z, cfg_lut_oflow_priority_rsc_z, cfg_lut_hybrid_priority_rsc_z,
      cfg_precision_rsc_z, chn_lut_out_rsc_z, chn_lut_out_rsc_vz, chn_lut_out_rsc_lz,
      chn_lut_in_rsci_oswt, chn_lut_in_rsci_oswt_unreg, chn_lut_out_rsci_oswt, chn_lut_out_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_lut_in_rsc_z;
  input chn_lut_in_rsc_vz;
  output chn_lut_in_rsc_lz;
  input [31:0] cfg_lut_le_start_rsc_z;
  input [31:0] cfg_lut_lo_start_rsc_z;
  input [7:0] cfg_lut_le_index_offset_rsc_z;
  input [7:0] cfg_lut_le_index_select_rsc_z;
  input [7:0] cfg_lut_lo_index_select_rsc_z;
  input cfg_lut_le_function_rsc_z;
  input cfg_lut_uflow_priority_rsc_z;
  input cfg_lut_oflow_priority_rsc_z;
  input cfg_lut_hybrid_priority_rsc_z;
  input [1:0] cfg_precision_rsc_z;
  output [323:0] chn_lut_out_rsc_z;
  input chn_lut_out_rsc_vz;
  output chn_lut_out_rsc_lz;
  input chn_lut_in_rsci_oswt;
  output chn_lut_in_rsci_oswt_unreg;
  input chn_lut_out_rsci_oswt;
  output chn_lut_out_rsci_oswt_unreg;


  // Interconnect Declarations
  wire core_wen;
  reg chn_lut_in_rsci_iswt0;
  wire chn_lut_in_rsci_bawt;
  wire chn_lut_in_rsci_wen_comp;
  reg chn_lut_in_rsci_ld_core_psct;
  wire [127:0] chn_lut_in_rsci_d_mxwt;
  wire core_wten;
  wire [31:0] cfg_lut_le_start_rsci_d;
  wire [31:0] cfg_lut_lo_start_rsci_d;
  wire [7:0] cfg_lut_le_index_offset_rsci_d;
  wire [7:0] cfg_lut_le_index_select_rsci_d;
  wire [7:0] cfg_lut_lo_index_select_rsci_d;
  wire cfg_lut_le_function_rsci_d;
  wire cfg_lut_uflow_priority_rsci_d;
  wire cfg_lut_oflow_priority_rsci_d;
  wire cfg_lut_hybrid_priority_rsci_d;
  wire [1:0] cfg_precision_rsci_d;
  reg chn_lut_out_rsci_iswt0;
  wire chn_lut_out_rsci_bawt;
  wire chn_lut_out_rsci_wen_comp;
  reg chn_lut_out_rsci_d_323;
  reg chn_lut_out_rsci_d_322;
  reg chn_lut_out_rsci_d_321;
  reg chn_lut_out_rsci_d_320;
  reg chn_lut_out_rsci_d_319;
  reg chn_lut_out_rsci_d_318;
  reg chn_lut_out_rsci_d_317;
  reg chn_lut_out_rsci_d_316;
  reg chn_lut_out_rsci_d_315;
  reg chn_lut_out_rsci_d_314;
  reg chn_lut_out_rsci_d_313;
  reg [5:0] chn_lut_out_rsci_d_312_307;
  reg chn_lut_out_rsci_d_306;
  reg chn_lut_out_rsci_d_305;
  reg chn_lut_out_rsci_d_304;
  reg [5:0] chn_lut_out_rsci_d_303_298;
  reg chn_lut_out_rsci_d_297;
  reg chn_lut_out_rsci_d_296;
  reg chn_lut_out_rsci_d_295;
  reg [5:0] chn_lut_out_rsci_d_294_289;
  reg chn_lut_out_rsci_d_288;
  reg chn_lut_out_rsci_d_287;
  reg chn_lut_out_rsci_d_286;
  reg [5:0] chn_lut_out_rsci_d_285_280;
  reg chn_lut_out_rsci_d_279;
  reg chn_lut_out_rsci_d_278;
  reg chn_lut_out_rsci_d_277;
  reg chn_lut_out_rsci_d_276;
  reg chn_lut_out_rsci_d_275;
  reg chn_lut_out_rsci_d_274;
  reg chn_lut_out_rsci_d_273;
  reg chn_lut_out_rsci_d_272;
  reg chn_lut_out_rsci_d_271;
  reg chn_lut_out_rsci_d_270;
  reg chn_lut_out_rsci_d_269;
  reg chn_lut_out_rsci_d_268;
  reg [127:0] chn_lut_out_rsci_d_267_140;
  reg [22:0] chn_lut_out_rsci_d_139_117;
  reg [11:0] chn_lut_out_rsci_d_116_105;
  reg [22:0] chn_lut_out_rsci_d_104_82;
  reg [11:0] chn_lut_out_rsci_d_81_70;
  reg [22:0] chn_lut_out_rsci_d_69_47;
  reg [11:0] chn_lut_out_rsci_d_46_35;
  reg [22:0] chn_lut_out_rsci_d_34_12;
  reg [11:0] chn_lut_out_rsci_d_11_0;
  wire [1:0] fsm_output;
  wire lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  wire IsNaN_8U_23U_3_nor_6_tmp;
  wire lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  wire IsNaN_8U_23U_3_nor_10_tmp;
  wire lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  wire IsNaN_8U_23U_3_nor_4_tmp;
  wire lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  wire IsNaN_8U_23U_3_nor_8_tmp;
  wire lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp;
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp;
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp;
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp;
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp;
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp;
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp;
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp;
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp;
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp;
  wire [7:0] FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp;
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp;
  wire [9:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [9:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [9:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [9:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [9:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [9:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [9:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  wire [9:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire [10:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  wire lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp;
  wire [8:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  wire lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp;
  wire lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp;
  wire [8:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  wire lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp;
  wire lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp;
  wire [8:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  wire lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp;
  wire lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp;
  wire [8:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  wire lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
  wire IsNaN_8U_23U_8_nor_2_tmp_1;
  wire IsNaN_8U_23U_4_nor_tmp;
  wire or_tmp_6;
  wire or_tmp_8;
  wire mux_tmp_4;
  wire mux_tmp_10;
  wire not_tmp_47;
  wire or_tmp_44;
  wire mux_tmp_35;
  wire or_tmp_63;
  wire and_tmp_5;
  wire and_tmp_6;
  wire or_tmp_101;
  wire nor_tmp_12;
  wire nor_tmp_14;
  wire or_tmp_124;
  wire mux_tmp_70;
  wire mux_tmp_72;
  wire or_tmp_129;
  wire mux_tmp_76;
  wire mux_tmp_78;
  wire nor_tmp_32;
  wire nor_tmp_34;
  wire mux_tmp_128;
  wire nand_tmp_4;
  wire and_tmp_14;
  wire nor_tmp_44;
  wire nor_tmp_46;
  wire and_tmp_19;
  wire nor_tmp_55;
  wire nor_tmp_57;
  wire mux_tmp_207;
  wire or_tmp_314;
  wire not_tmp_209;
  wire mux_tmp_220;
  wire or_tmp_331;
  wire and_tmp_27;
  wire not_tmp_222;
  wire or_tmp_363;
  wire not_tmp_235;
  wire or_tmp_378;
  wire or_tmp_380;
  wire or_tmp_395;
  wire or_tmp_397;
  wire not_tmp_248;
  wire or_tmp_427;
  wire or_tmp_428;
  wire mux_tmp_265;
  wire or_tmp_447;
  wire mux_tmp_270;
  wire or_tmp_456;
  wire mux_tmp_279;
  wire mux_tmp_281;
  wire or_tmp_478;
  wire not_tmp_276;
  wire mux_tmp_292;
  wire or_tmp_505;
  wire or_tmp_522;
  wire mux_tmp_301;
  wire or_tmp_547;
  wire or_tmp_573;
  wire or_tmp_598;
  wire or_tmp_623;
  wire not_tmp_334;
  wire nor_tmp_112;
  wire mux_tmp_475;
  wire not_tmp_394;
  wire not_tmp_412;
  wire not_tmp_418;
  wire not_tmp_422;
  wire mux_tmp_595;
  wire mux_tmp_596;
  wire or_tmp_843;
  wire mux_tmp_617;
  wire mux_tmp_618;
  wire mux_tmp_643;
  wire and_tmp_59;
  wire and_tmp_61;
  wire mux_tmp_655;
  wire and_tmp_69;
  wire mux_tmp_704;
  wire and_tmp_83;
  wire or_tmp_976;
  wire or_tmp_980;
  wire or_tmp_993;
  wire and_tmp_92;
  wire nor_tmp_238;
  wire and_tmp_97;
  wire or_tmp_1043;
  wire and_tmp_98;
  wire and_tmp_103;
  wire nor_tmp_260;
  wire nand_tmp_22;
  wire and_tmp_108;
  wire and_tmp_113;
  wire nor_tmp_281;
  wire or_tmp_1181;
  wire and_tmp_119;
  wire and_tmp_124;
  wire and_tmp_130;
  wire or_tmp_1250;
  wire and_tmp_131;
  wire mux_tmp_978;
  wire or_tmp_1360;
  wire not_tmp_800;
  wire or_tmp_1450;
  wire mux_tmp_1101;
  wire mux_tmp_1104;
  wire and_tmp_178;
  wire and_dcpl_54;
  wire and_dcpl_59;
  wire and_dcpl_63;
  wire and_dcpl_67;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_74;
  wire or_tmp_1490;
  wire and_dcpl_98;
  wire and_dcpl_148;
  wire or_dcpl_51;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire or_dcpl_57;
  wire mux_tmp_1130;
  wire or_tmp_1513;
  wire mux_tmp_1136;
  wire mux_tmp_1143;
  wire or_tmp_1523;
  wire mux_tmp_1149;
  wire mux_tmp_1156;
  wire or_tmp_1534;
  wire mux_tmp_1162;
  wire mux_tmp_1169;
  wire or_tmp_1545;
  wire mux_tmp_1175;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire and_dcpl_280;
  wire and_dcpl_284;
  wire and_dcpl_288;
  wire and_dcpl_292;
  wire and_dcpl_296;
  wire and_dcpl_300;
  wire and_dcpl_304;
  wire and_dcpl_308;
  wire and_dcpl_309;
  wire and_dcpl_314;
  wire and_dcpl_315;
  wire and_dcpl_316;
  wire and_dcpl_351;
  wire and_dcpl_364;
  wire and_dcpl_403;
  wire and_dcpl_405;
  wire or_tmp_1628;
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2;
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1;
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1;
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_sva_1;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg main_stage_v_5;
  reg IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  reg IsNaN_8U_23U_8_land_lpi_1_dfm_5;
  reg lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_8_land_3_lpi_1_dfm_4;
  reg IsNaN_8U_23U_8_land_3_lpi_1_dfm_5;
  reg lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_3_lpi_1_dfm_5;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  reg IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  reg lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_2_lpi_1_dfm_5;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_8_land_1_lpi_1_dfm_7;
  reg lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  reg IsNaN_8U_23U_4_land_1_lpi_1_dfm_4;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  reg lut_lookup_4_if_else_slc_32_svs_5;
  reg lut_lookup_4_if_else_slc_32_svs_6;
  reg lut_lookup_4_if_else_slc_32_svs_7;
  reg lut_lookup_4_if_else_slc_32_svs_8;
  reg lut_lookup_3_if_else_slc_32_svs_5;
  reg lut_lookup_3_if_else_slc_32_svs_6;
  reg lut_lookup_3_if_else_slc_32_svs_7;
  reg lut_lookup_3_if_else_slc_32_svs_8;
  reg lut_lookup_2_if_else_slc_32_svs_5;
  reg lut_lookup_2_if_else_slc_32_svs_6;
  reg lut_lookup_2_if_else_slc_32_svs_7;
  reg lut_lookup_2_if_else_slc_32_svs_8;
  reg lut_lookup_1_if_else_slc_32_svs_5;
  reg lut_lookup_1_if_else_slc_32_svs_6;
  reg lut_lookup_1_if_else_slc_32_svs_7;
  reg lut_lookup_1_if_else_slc_32_svs_8;
  reg lut_lookup_else_unequal_tmp_12;
  reg lut_lookup_else_unequal_tmp_13;
  reg lut_lookup_else_unequal_tmp_18;
  reg [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_11;
  reg [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_12;
  reg [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_13;
  reg [34:0] lut_lookup_lo_fraction_lpi_1_dfm_9;
  reg lut_lookup_else_1_slc_32_mdf_sva_5;
  reg lut_lookup_else_1_slc_32_mdf_sva_6;
  reg lut_lookup_else_1_slc_32_mdf_sva_7;
  reg lut_lookup_else_1_slc_32_mdf_sva_8;
  reg [34:0] lut_lookup_if_1_else_lo_fra_sva_4;
  reg lut_lookup_if_1_lor_1_lpi_1_dfm_4;
  reg lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_sva_3;
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_25;
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_26;
  reg [34:0] lut_lookup_le_fraction_lpi_1_dfm_21;
  reg lut_lookup_else_else_else_asn_mdf_sva_3;
  reg lut_lookup_else_else_else_asn_mdf_sva_4;
  reg lut_lookup_else_else_slc_32_mdf_sva_7;
  reg lut_lookup_else_else_slc_32_mdf_sva_8;
  reg [34:0] lut_lookup_else_if_else_le_fra_sva_4;
  reg lut_lookup_else_if_lor_1_lpi_1_dfm_5;
  reg lut_lookup_else_if_lor_1_lpi_1_dfm_6;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_sva_3;
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_27;
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_28;
  reg [34:0] lut_lookup_le_fraction_lpi_1_dfm_22;
  reg lut_lookup_if_else_else_else_asn_mdf_sva_2;
  reg lut_lookup_if_else_else_slc_10_mdf_sva_3;
  reg lut_lookup_if_else_else_slc_10_mdf_sva_4;
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_29;
  reg [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11;
  reg [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12;
  reg [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13;
  reg [34:0] lut_lookup_lo_fraction_3_lpi_1_dfm_9;
  reg lut_lookup_else_1_slc_32_mdf_3_sva_5;
  reg lut_lookup_else_1_slc_32_mdf_3_sva_6;
  reg lut_lookup_else_1_slc_32_mdf_3_sva_7;
  reg lut_lookup_else_1_slc_32_mdf_3_sva_8;
  reg [34:0] lut_lookup_if_1_else_lo_fra_3_sva_4;
  reg lut_lookup_if_1_lor_7_lpi_1_dfm_4;
  reg lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_3_sva_3;
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25;
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26;
  reg [34:0] lut_lookup_le_fraction_3_lpi_1_dfm_21;
  reg lut_lookup_else_else_else_asn_mdf_3_sva_3;
  reg lut_lookup_else_else_else_asn_mdf_3_sva_4;
  reg lut_lookup_else_else_slc_32_mdf_3_sva_7;
  reg lut_lookup_else_else_slc_32_mdf_3_sva_8;
  reg [34:0] lut_lookup_else_if_else_le_fra_3_sva_4;
  reg lut_lookup_else_if_lor_7_lpi_1_dfm_5;
  reg lut_lookup_else_if_lor_7_lpi_1_dfm_6;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_3_sva_3;
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27;
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28;
  reg [34:0] lut_lookup_le_fraction_3_lpi_1_dfm_22;
  reg lut_lookup_if_else_else_else_asn_mdf_3_sva_2;
  reg lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  reg lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29;
  reg [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11;
  reg [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12;
  reg [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13;
  reg [34:0] lut_lookup_lo_fraction_2_lpi_1_dfm_9;
  reg lut_lookup_else_1_slc_32_mdf_2_sva_5;
  reg lut_lookup_else_1_slc_32_mdf_2_sva_6;
  reg lut_lookup_else_1_slc_32_mdf_2_sva_7;
  reg lut_lookup_else_1_slc_32_mdf_2_sva_8;
  reg [34:0] lut_lookup_if_1_else_lo_fra_2_sva_4;
  reg lut_lookup_if_1_lor_6_lpi_1_dfm_4;
  reg lut_lookup_if_1_lor_6_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_2_sva_3;
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25;
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26;
  reg [34:0] lut_lookup_le_fraction_2_lpi_1_dfm_21;
  reg lut_lookup_else_else_else_asn_mdf_2_sva_3;
  reg lut_lookup_else_else_else_asn_mdf_2_sva_4;
  reg lut_lookup_else_else_slc_32_mdf_2_sva_7;
  reg lut_lookup_else_else_slc_32_mdf_2_sva_8;
  reg [34:0] lut_lookup_else_if_else_le_fra_2_sva_4;
  reg lut_lookup_else_if_lor_6_lpi_1_dfm_5;
  reg lut_lookup_else_if_lor_6_lpi_1_dfm_6;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_2_sva_3;
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27;
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28;
  reg [34:0] lut_lookup_le_fraction_2_lpi_1_dfm_22;
  reg lut_lookup_if_else_else_else_asn_mdf_2_sva_2;
  reg lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  reg lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29;
  reg [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11;
  reg [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12;
  reg [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13;
  reg [34:0] lut_lookup_lo_fraction_1_lpi_1_dfm_9;
  reg lut_lookup_else_1_slc_32_mdf_1_sva_5;
  reg lut_lookup_else_1_slc_32_mdf_1_sva_6;
  reg lut_lookup_else_1_slc_32_mdf_1_sva_7;
  reg lut_lookup_else_1_slc_32_mdf_1_sva_8;
  reg [34:0] lut_lookup_if_1_else_lo_fra_1_sva_4;
  reg lut_lookup_if_1_lor_5_lpi_1_dfm_4;
  reg lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_1_sva_3;
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25;
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26;
  reg [34:0] lut_lookup_le_fraction_1_lpi_1_dfm_21;
  reg lut_lookup_else_else_else_asn_mdf_1_sva_3;
  reg lut_lookup_else_else_else_asn_mdf_1_sva_4;
  reg lut_lookup_else_else_slc_32_mdf_1_sva_7;
  reg lut_lookup_else_else_slc_32_mdf_1_sva_8;
  reg [34:0] lut_lookup_else_if_else_le_fra_1_sva_4;
  reg lut_lookup_else_if_lor_5_lpi_1_dfm_5;
  reg lut_lookup_else_if_lor_5_lpi_1_dfm_6;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_1_sva_3;
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3;
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27;
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28;
  reg [34:0] lut_lookup_le_fraction_1_lpi_1_dfm_22;
  reg lut_lookup_if_else_else_else_asn_mdf_1_sva_2;
  reg lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  reg lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29;
  reg [31:0] cfg_lut_le_start_1_sva_41;
  reg [31:0] cfg_lut_lo_start_1_sva_41;
  reg [7:0] cfg_lut_le_index_offset_1_sva_4;
  reg [7:0] cfg_lut_le_index_offset_1_sva_5;
  reg [7:0] cfg_lut_le_index_offset_1_sva_6;
  reg [7:0] cfg_lut_le_index_offset_1_sva_7;
  reg [7:0] cfg_lut_le_index_select_1_sva_4;
  reg [7:0] cfg_lut_le_index_select_1_sva_5;
  reg [7:0] cfg_lut_le_index_select_1_sva_6;
  reg [7:0] cfg_lut_lo_index_select_1_sva_4;
  reg [7:0] cfg_lut_lo_index_select_1_sva_5;
  reg [7:0] cfg_lut_lo_index_select_1_sva_6;
  reg cfg_lut_le_function_1_sva_10;
  reg cfg_lut_uflow_priority_1_sva_6;
  reg cfg_lut_uflow_priority_1_sva_7;
  reg cfg_lut_uflow_priority_1_sva_8;
  reg cfg_lut_uflow_priority_1_sva_9;
  reg cfg_lut_uflow_priority_1_sva_10;
  reg cfg_lut_oflow_priority_1_sva_6;
  reg cfg_lut_oflow_priority_1_sva_7;
  reg cfg_lut_oflow_priority_1_sva_8;
  reg cfg_lut_oflow_priority_1_sva_9;
  reg cfg_lut_oflow_priority_1_sva_10;
  reg cfg_lut_hybrid_priority_1_sva_6;
  reg cfg_lut_hybrid_priority_1_sva_7;
  reg cfg_lut_hybrid_priority_1_sva_8;
  reg cfg_lut_hybrid_priority_1_sva_9;
  reg cfg_lut_hybrid_priority_1_sva_10;
  reg [1:0] cfg_precision_1_sva_8;
  reg [127:0] lut_in_data_sva_154;
  reg [127:0] lut_in_data_sva_155;
  reg [127:0] lut_in_data_sva_156;
  reg [127:0] lut_in_data_sva_157;
  reg [127:0] lut_in_data_sva_158;
  reg FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5;
  reg FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  reg FpMantRNE_49U_24U_1_else_carry_1_sva_2;
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2;
  reg IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_6_land_1_lpi_1_dfm_7;
  reg [31:0] lut_lookup_else_else_else_le_index_u_1_sva_3;
  reg [31:0] lut_lookup_else_else_else_le_index_u_1_sva_4;
  reg lut_lookup_le_uflow_1_lpi_1_dfm_6;
  reg lut_lookup_unequal_tmp_13;
  reg FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12;
  reg FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  reg FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  reg lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2;
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  reg [22:0] FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2;
  reg IsNaN_8U_23U_10_land_1_lpi_1_dfm_5;
  reg IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  reg [31:0] lut_lookup_else_1_lo_index_u_1_sva_3;
  wire [32:0] nl_lut_lookup_else_1_lo_index_u_1_sva_3;
  reg [31:0] lut_lookup_else_1_lo_index_u_1_sva_4;
  reg lut_lookup_lo_uflow_1_lpi_1_dfm_3;
  reg lut_lookup_lo_uflow_1_lpi_1_dfm_4;
  reg lut_lookup_1_and_svs_2;
  reg FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5;
  reg FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  reg FpMantRNE_49U_24U_1_else_carry_2_sva_2;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2;
  reg IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_6_land_2_lpi_1_dfm_7;
  reg [31:0] lut_lookup_else_else_else_le_index_u_2_sva_3;
  reg [31:0] lut_lookup_else_else_else_le_index_u_2_sva_4;
  reg lut_lookup_le_uflow_2_lpi_1_dfm_6;
  reg FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12;
  reg FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  reg FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  reg lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  reg [22:0] FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2;
  reg IsNaN_8U_23U_10_land_2_lpi_1_dfm_5;
  reg IsNaN_8U_23U_10_land_2_lpi_1_dfm_6;
  reg [31:0] lut_lookup_else_1_lo_index_u_2_sva_3;
  wire [32:0] nl_lut_lookup_else_1_lo_index_u_2_sva_3;
  reg [31:0] lut_lookup_else_1_lo_index_u_2_sva_4;
  reg lut_lookup_lo_uflow_2_lpi_1_dfm_3;
  reg lut_lookup_lo_uflow_2_lpi_1_dfm_4;
  reg lut_lookup_2_and_svs_2;
  reg FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5;
  reg FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  reg FpMantRNE_49U_24U_1_else_carry_3_sva_2;
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2;
  reg IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  reg IsNaN_8U_23U_6_land_3_lpi_1_dfm_7;
  reg [31:0] lut_lookup_else_else_else_le_index_u_3_sva_3;
  reg [31:0] lut_lookup_else_else_else_le_index_u_3_sva_4;
  reg lut_lookup_le_uflow_3_lpi_1_dfm_6;
  reg FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12;
  reg FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  reg FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  reg lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2;
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  reg [22:0] FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2;
  reg IsNaN_8U_23U_10_land_3_lpi_1_dfm_5;
  reg IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  reg [31:0] lut_lookup_else_1_lo_index_u_3_sva_3;
  wire [32:0] nl_lut_lookup_else_1_lo_index_u_3_sva_3;
  reg [31:0] lut_lookup_else_1_lo_index_u_3_sva_4;
  reg lut_lookup_lo_uflow_3_lpi_1_dfm_3;
  reg lut_lookup_lo_uflow_3_lpi_1_dfm_4;
  reg lut_lookup_3_and_svs_2;
  reg FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_1_qr_lpi_1_dfm_5;
  reg FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  reg FpMantRNE_49U_24U_1_else_carry_sva_2;
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2;
  reg IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_6_land_lpi_1_dfm_7;
  reg [31:0] lut_lookup_else_else_else_le_index_u_sva_3;
  reg [31:0] lut_lookup_else_else_else_le_index_u_sva_4;
  reg lut_lookup_le_uflow_lpi_1_dfm_6;
  reg FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_lpi_1_dfm_4;
  reg [7:0] FpAdd_8U_23U_2_qr_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12;
  reg FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  reg FpMantRNE_49U_24U_2_else_carry_sva_2;
  reg lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2;
  reg IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  reg [22:0] FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5;
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2;
  reg IsNaN_8U_23U_10_land_lpi_1_dfm_5;
  reg IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  reg [31:0] lut_lookup_else_1_lo_index_u_sva_3;
  wire [32:0] nl_lut_lookup_else_1_lo_index_u_sva_3;
  reg [31:0] lut_lookup_else_1_lo_index_u_sva_4;
  reg lut_lookup_lo_uflow_lpi_1_dfm_3;
  reg lut_lookup_lo_uflow_lpi_1_dfm_4;
  reg lut_lookup_4_and_svs_2;
  reg [1:0] lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  reg [5:0] lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  reg lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  reg IsNaN_8U_23U_4_nor_itm_2;
  reg IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2;
  reg [22:0] lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  reg FpAdd_8U_23U_1_mux_1_itm_2;
  reg FpAdd_8U_23U_1_mux_13_itm_3;
  reg FpAdd_8U_23U_1_mux_13_itm_4;
  reg [7:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  reg lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  reg [31:0] lut_lookup_1_else_else_else_else_le_data_f_and_itm_2;
  reg lut_lookup_else_mux_itm_2;
  reg lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2;
  reg lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  reg [22:0] lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  reg FpAdd_8U_23U_2_mux_1_itm_2;
  reg FpAdd_8U_23U_2_mux_13_itm_1;
  reg FpAdd_8U_23U_2_mux_13_itm_3;
  reg [7:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  wire [8:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  reg lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  reg [31:0] lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2;
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  reg lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2;
  reg [1:0] lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  reg [5:0] lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  reg lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  reg [22:0] lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  reg FpAdd_8U_23U_1_mux_17_itm_2;
  reg FpAdd_8U_23U_1_mux_29_itm_3;
  reg FpAdd_8U_23U_1_mux_29_itm_4;
  reg [7:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  reg lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  reg [31:0] lut_lookup_2_else_else_else_else_le_data_f_and_itm_2;
  reg lut_lookup_else_mux_43_itm_2;
  reg lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2;
  reg lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  reg [22:0] lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  reg FpAdd_8U_23U_2_mux_17_itm_2;
  reg FpAdd_8U_23U_2_mux_29_itm_1;
  reg FpAdd_8U_23U_2_mux_29_itm_3;
  reg [7:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  wire [8:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  reg lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  reg [31:0] lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2;
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  reg lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2;
  reg [1:0] lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  reg [5:0] lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  reg lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  reg [22:0] lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  reg FpAdd_8U_23U_1_mux_33_itm_2;
  reg FpAdd_8U_23U_1_mux_45_itm_3;
  reg FpAdd_8U_23U_1_mux_45_itm_4;
  reg [7:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  reg lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  reg [31:0] lut_lookup_3_else_else_else_else_le_data_f_and_itm_2;
  reg lut_lookup_else_mux_86_itm_2;
  reg lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2;
  reg lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  reg IsNaN_8U_23U_8_nor_2_itm_2;
  reg IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2;
  reg [22:0] lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  reg FpAdd_8U_23U_2_mux_33_itm_2;
  reg FpAdd_8U_23U_2_mux_45_itm_1;
  reg FpAdd_8U_23U_2_mux_45_itm_3;
  reg [7:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  wire [8:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  reg lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  reg [31:0] lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2;
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  reg lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2;
  reg [1:0] lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  reg [5:0] lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  reg lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  reg IsNaN_8U_23U_4_nor_3_itm_2;
  reg IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2;
  reg [22:0] lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  reg FpAdd_8U_23U_1_mux_49_itm_2;
  reg FpAdd_8U_23U_1_mux_61_itm_3;
  reg FpAdd_8U_23U_1_mux_61_itm_4;
  reg [7:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  reg lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  reg [31:0] lut_lookup_4_else_else_else_else_le_data_f_and_itm_2;
  reg lut_lookup_else_mux_129_itm_2;
  reg lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2;
  reg lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  reg lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2;
  reg IsNaN_8U_23U_8_nor_3_itm_2;
  reg IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2;
  reg [22:0] lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  reg FpAdd_8U_23U_2_mux_49_itm_2;
  reg FpAdd_8U_23U_2_mux_61_itm_1;
  reg FpAdd_8U_23U_2_mux_61_itm_3;
  reg [7:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  wire [8:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  reg lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  reg [31:0] lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2;
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  reg lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2;
  reg lut_lookup_else_2_else_else_if_mux_26_itm_1;
  reg lut_lookup_else_2_else_else_if_mux_19_itm_1;
  reg lut_lookup_else_2_else_else_if_mux_12_itm_1;
  reg lut_lookup_else_2_else_else_if_mux_5_itm_1;
  reg [1:0] cfg_precision_1_sva_st_70;
  reg [1:0] cfg_precision_1_sva_st_71;
  reg lut_lookup_1_if_else_slc_32_svs_st_5;
  reg lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3;
  reg lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6;
  reg [1:0] cfg_precision_1_sva_st_72;
  reg lut_lookup_else_if_lor_5_lpi_1_dfm_st_3;
  reg lut_lookup_else_else_else_asn_mdf_1_sva_st_3;
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6;
  reg lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  reg lut_lookup_2_if_else_slc_32_svs_st_5;
  reg lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3;
  reg lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6;
  reg lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  reg lut_lookup_else_else_else_asn_mdf_2_sva_st_3;
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6;
  reg lut_lookup_if_1_lor_6_lpi_1_dfm_st_4;
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  reg lut_lookup_3_if_else_slc_32_svs_st_5;
  reg lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3;
  reg lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6;
  reg lut_lookup_else_if_lor_7_lpi_1_dfm_st_3;
  reg lut_lookup_else_else_else_asn_mdf_3_sva_st_3;
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6;
  reg lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  reg cfg_lut_le_function_1_sva_st_41;
  reg cfg_lut_le_function_1_sva_st_42;
  reg lut_lookup_4_if_else_slc_32_svs_st_5;
  reg lut_lookup_if_else_else_slc_10_mdf_sva_st_3;
  reg lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_st_6;
  reg lut_lookup_else_if_lor_1_lpi_1_dfm_st_3;
  reg lut_lookup_else_else_else_asn_mdf_sva_st_3;
  reg IsNaN_8U_23U_7_land_lpi_1_dfm_st_6;
  reg [1:0] cfg_precision_1_sva_st_107;
  reg lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  reg [22:0] lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1;
  reg [22:0] lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1;
  reg [22:0] lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1;
  reg [22:0] lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1;
  reg [30:0] cfg_lut_le_start_1_sva_2_30_0_1;
  reg [30:0] cfg_lut_le_start_1_sva_3_30_0_1;
  reg [30:0] cfg_lut_lo_start_1_sva_2_30_0_1;
  reg [30:0] cfg_lut_lo_start_1_sva_3_30_0_1;
  reg [30:0] lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1;
  reg [30:0] lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1;
  reg [30:0] lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1;
  reg [30:0] lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1;
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1;
  wire main_stage_en_1;
  wire FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  wire FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  wire FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  wire FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  wire lut_lookup_or_3_tmp;
  wire lut_lookup_or_7_tmp;
  wire lut_lookup_or_11_tmp;
  wire lut_lookup_or_15_tmp;
  wire lut_lookup_le_miss_1_sva;
  wire lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  wire lut_lookup_1_else_2_and_svs;
  wire lut_lookup_le_miss_2_sva;
  wire lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  wire lut_lookup_2_else_2_and_svs;
  wire lut_lookup_le_miss_3_sva;
  wire lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  wire lut_lookup_3_else_2_and_svs;
  wire lut_lookup_le_miss_sva;
  wire lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  wire lut_lookup_4_else_2_and_svs;
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse;
  wire lut_lookup_lo_miss_sva;
  wire lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  wire lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0;
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse;
  wire lut_lookup_lo_miss_3_sva;
  wire lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  wire lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0;
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse;
  wire lut_lookup_lo_miss_2_sva;
  wire lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  wire lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0;
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse;
  wire lut_lookup_lo_miss_1_sva;
  wire lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  wire lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0;
  wire IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0;
  wire FpAdd_8U_23U_1_and_3_tmp;
  wire FpAdd_8U_23U_1_and_2_tmp;
  wire FpAdd_8U_23U_1_and_1_tmp;
  wire lut_lookup_if_mux_123_mx0w1;
  wire lut_lookup_if_mux_82_mx0w1;
  wire lut_lookup_if_mux_41_mx0w1;
  wire lut_lookup_if_mux_mx0w1;
  wire [8:0] lut_lookup_else_if_else_le_int_lpi_1_dfm_1;
  wire [8:0] lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1;
  wire [8:0] lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1;
  wire [8:0] lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1;
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_sva;
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_sva;
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_3_sva;
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_3_sva;
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_2_sva;
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_2_sva;
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_1_sva;
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_1_sva;
  wire [22:0] FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0;
  wire [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_7;
  wire [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7;
  wire [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7;
  wire and_597_m1c;
  wire and_590_m1c;
  wire and_592_m1c;
  wire and_582_m1c;
  wire and_577_m1c;
  wire and_572_m1c;
  wire and_567_m1c;
  wire and_562_m1c;
  wire and_553_m1c;
  wire and_555_m1c;
  wire and_375_m1c;
  wire and_355_m1c;
  wire chn_lut_out_and_cse;
  wire chn_lut_out_and_13_cse;
  wire chn_lut_out_and_14_cse;
  wire chn_lut_out_and_15_cse;
  wire chn_lut_out_and_16_cse;
  wire nor_13_cse;
  wire nor_31_cse;
  wire nor_42_cse;
  wire nor_54_cse;
  wire and_854_cse;
  wire and_846_cse;
  wire and_82_cse;
  wire and_839_cse;
  wire and_835_cse;
  wire lut_lookup_else_mux_180_cse;
  wire lut_lookup_else_mux_182_cse;
  wire lut_lookup_else_mux_184_cse;
  wire lut_lookup_else_mux_186_cse;
  wire and_465_cse;
  wire and_466_cse;
  wire or_1853_cse;
  reg reg_chn_lut_out_rsci_ld_core_psct_cse;
  wire or_26_cse;
  wire nor_648_cse;
  wire or_1857_cse;
  wire or_978_cse;
  wire nor_612_cse;
  wire and_814_cse;
  wire and_811_cse;
  wire or_66_cse;
  wire and_795_cse;
  wire and_789_cse;
  wire and_787_cse;
  wire and_784_cse;
  wire and_794_cse;
  wire and_780_cse;
  wire or_969_cse;
  wire nor_469_cse;
  wire nor_482_cse;
  wire lut_lookup_and_138_cse;
  wire lut_lookup_and_139_cse;
  wire lut_lookup_and_136_cse;
  wire lut_lookup_and_137_cse;
  wire lut_lookup_and_134_cse;
  wire lut_lookup_and_135_cse;
  wire lut_lookup_and_132_cse;
  wire lut_lookup_and_133_cse;
  wire or_1689_cse;
  wire and_850_cse;
  wire and_848_cse;
  wire nor_610_cse;
  wire nor_526_cse;
  wire lut_lookup_if_else_lut_lookup_if_else_or_cse;
  wire lut_lookup_if_else_lut_lookup_if_else_or_1_cse;
  wire lut_lookup_if_else_lut_lookup_if_else_or_2_cse;
  wire lut_lookup_if_else_lut_lookup_if_else_or_3_cse;
  wire or_1202_cse;
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse;
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse;
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse;
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse;
  wire or_1495_cse;
  wire lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1;
  wire IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
  wire [8:0] lut_lookup_else_else_else_else_mux1h_rgt;
  wire [30:0] IntLog2_32U_IntLog2_32U_mux_rgt;
  wire [8:0] lut_lookup_else_else_else_else_mux1h_1_rgt;
  wire [30:0] IntLog2_32U_IntLog2_32U_mux_1_rgt;
  wire [8:0] lut_lookup_else_else_else_else_mux1h_2_rgt;
  wire [30:0] IntLog2_32U_IntLog2_32U_mux_2_rgt;
  wire [8:0] lut_lookup_else_else_else_else_mux1h_3_rgt;
  reg reg_lut_lookup_1_else_else_else_else_acc_reg;
  reg reg_lut_lookup_1_else_else_else_else_acc_1_reg;
  reg [2:0] reg_lut_lookup_1_else_else_else_else_acc_2_reg;
  reg [3:0] reg_lut_lookup_1_else_else_else_else_acc_3_reg;
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg;
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg;
  reg reg_lut_lookup_2_else_else_else_else_acc_reg;
  reg reg_lut_lookup_2_else_else_else_else_acc_1_reg;
  reg [2:0] reg_lut_lookup_2_else_else_else_else_acc_2_reg;
  reg [3:0] reg_lut_lookup_2_else_else_else_else_acc_3_reg;
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg;
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg;
  reg reg_lut_lookup_3_else_else_else_else_acc_reg;
  reg reg_lut_lookup_3_else_else_else_else_acc_1_reg;
  reg [2:0] reg_lut_lookup_3_else_else_else_else_acc_2_reg;
  reg [3:0] reg_lut_lookup_3_else_else_else_else_acc_3_reg;
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_reg;
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1;
  reg reg_lut_lookup_4_else_else_else_else_acc_reg;
  reg reg_lut_lookup_4_else_else_else_else_acc_1_reg;
  reg [2:0] reg_lut_lookup_4_else_else_else_else_acc_2_reg;
  reg [3:0] reg_lut_lookup_4_else_else_else_else_acc_3_reg;
  wire mux_789_cse;
  wire mux_845_cse;
  wire mux_900_cse;
  wire mux_959_cse;
  wire [7:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0;
  wire [8:0] nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0;
  wire [22:0] FpAdd_8U_23U_asn_45_mx0w1;
  wire [22:0] FpAdd_8U_23U_asn_40_mx0w1;
  wire [22:0] FpAdd_8U_23U_asn_35_mx0w1;
  wire mux_755_cse;
  wire and_896_cse;
  wire nor_588_cse;
  wire nor_564_cse;
  wire and_905_cse;
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_1_sva;
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_1_sva;
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_2_sva;
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_2_sva;
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_3_sva;
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_3_sva;
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_sva;
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_sva;
  wire and_dcpl_540;
  wire and_284_rgt;
  wire and_286_rgt;
  wire and_288_rgt;
  wire and_290_rgt;
  wire and_292_rgt;
  wire and_300_rgt;
  wire and_302_rgt;
  wire and_304_rgt;
  wire and_306_rgt;
  wire and_308_rgt;
  wire and_316_rgt;
  wire and_318_rgt;
  wire and_320_rgt;
  wire and_322_rgt;
  wire and_324_rgt;
  wire and_330_rgt;
  wire and_332_rgt;
  wire and_334_rgt;
  wire and_336_rgt;
  wire and_338_rgt;
  wire and_344_rgt;
  wire and_347_rgt;
  wire or_tmp_1663;
  wire and_dcpl_576;
  wire or_tmp_1671;
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt;
  wire FpAdd_8U_23U_2_and_4_rgt;
  wire FpAdd_8U_23U_2_and_5_rgt;
  wire and_364_rgt;
  wire or_tmp_1674;
  wire or_tmp_1678;
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt;
  wire FpAdd_8U_23U_2_and_10_rgt;
  wire FpAdd_8U_23U_2_and_11_rgt;
  wire or_tmp_1684;
  wire or_tmp_1692;
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt;
  wire FpAdd_8U_23U_2_and_16_rgt;
  wire FpAdd_8U_23U_2_and_17_rgt;
  wire or_tmp_1697;
  wire or_tmp_1705;
  wire or_tmp_1707;
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt;
  wire FpAdd_8U_23U_2_and_22_rgt;
  wire FpAdd_8U_23U_2_and_23_rgt;
  wire and_428_rgt;
  wire and_430_rgt;
  wire and_524_rgt;
  wire and_525_rgt;
  wire and_527_rgt;
  wire and_529_rgt;
  wire and_551_rgt;
  wire lut_lookup_or_17_rgt;
  wire lut_lookup_or_18_rgt;
  wire and_559_rgt;
  wire lut_lookup_and_126_rgt;
  wire lut_lookup_and_127_rgt;
  wire and_564_rgt;
  wire and_566_rgt;
  wire lut_lookup_and_124_rgt;
  wire lut_lookup_and_125_rgt;
  wire and_570_rgt;
  wire lut_lookup_and_122_rgt;
  wire lut_lookup_and_123_rgt;
  wire and_574_rgt;
  wire and_576_rgt;
  wire lut_lookup_and_120_rgt;
  wire lut_lookup_and_121_rgt;
  wire and_580_rgt;
  wire lut_lookup_and_118_rgt;
  wire lut_lookup_and_119_rgt;
  wire and_586_rgt;
  wire and_588_rgt;
  wire lut_lookup_or_rgt;
  wire lut_lookup_or_16_rgt;
  wire and_595_rgt;
  wire lut_lookup_and_112_rgt;
  wire lut_lookup_and_113_rgt;
  wire and_604_rgt;
  wire and_606_rgt;
  wire and_dcpl_648;
  wire and_653_rgt;
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp;
  wire or_tmp_1716;
  wire and_661_rgt;
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp;
  wire or_tmp_1720;
  wire and_668_rgt;
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp;
  wire and_676_rgt;
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp;
  wire and_679_rgt;
  wire [7:0] FpAdd_8U_23U_1_mux1h_1_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm;
  wire [7:0] FpAdd_8U_23U_1_mux1h_3_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm;
  wire [7:0] FpAdd_8U_23U_1_mux1h_5_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm;
  wire [7:0] FpAdd_8U_23U_1_mux1h_7_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm;
  reg reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  reg [1:0] reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm;
  reg reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  reg [1:0] reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm;
  reg reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  reg [1:0] reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm;
  reg reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  reg [1:0] reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm;
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm;
  wire [34:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  wire [255:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  wire [34:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  wire [255:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  wire [34:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  wire [255:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  wire [34:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  wire [255:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  wire [34:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  wire [255:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  wire [34:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  wire [255:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  wire [34:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  wire [255:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  wire [34:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  wire [255:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  wire [34:0] lut_lookup_1_if_else_else_else_else_if_lshift_itm;
  wire [34:0] lut_lookup_1_if_else_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_1_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_1_else_1_else_else_rshift_itm;
  wire [34:0] lut_lookup_2_if_else_else_else_else_if_lshift_itm;
  wire [34:0] lut_lookup_2_if_else_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_2_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_2_else_1_else_else_rshift_itm;
  wire [34:0] lut_lookup_3_if_else_else_else_else_if_lshift_itm;
  wire [34:0] lut_lookup_3_if_else_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_3_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_3_else_1_else_else_rshift_itm;
  wire [34:0] lut_lookup_4_if_else_else_else_else_if_lshift_itm;
  wire [34:0] lut_lookup_4_if_else_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_4_else_else_else_else_rshift_itm;
  wire [34:0] lut_lookup_4_else_1_else_else_rshift_itm;
  wire [30:0] IntLog2_32U_mux1h_1_itm;
  wire [30:0] lut_lookup_1_IntLog2_32U_lshift_itm;
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm;
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm;
  wire [8:0] lut_lookup_else_1_else_else_mux1h_1_itm;
  reg reg_lut_lookup_1_else_1_else_else_acc_itm;
  reg [7:0] reg_lut_lookup_1_else_1_else_else_acc_1_itm;
  wire [30:0] lut_lookup_2_IntLog2_32U_lshift_itm;
  reg reg_lut_lookup_2_else_1_else_else_acc_itm;
  reg [7:0] reg_lut_lookup_2_else_1_else_else_acc_1_itm;
  wire [30:0] lut_lookup_3_IntLog2_32U_lshift_itm;
  reg reg_lut_lookup_3_else_1_else_else_acc_itm;
  reg [7:0] reg_lut_lookup_3_else_1_else_else_acc_1_itm;
  wire [30:0] lut_lookup_4_IntLog2_32U_lshift_itm;
  reg reg_lut_lookup_4_else_1_else_else_acc_itm;
  reg [7:0] reg_lut_lookup_4_else_1_else_else_acc_1_itm;
  wire [48:0] lut_lookup_1_FpNormalize_8U_49U_else_lshift_itm;
  wire [286:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_itm;
  wire [286:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_2_FpNormalize_8U_49U_else_lshift_itm;
  wire [286:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_itm;
  wire [286:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_3_FpNormalize_8U_49U_else_lshift_itm;
  wire [286:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_itm;
  wire [286:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_4_FpNormalize_8U_49U_else_lshift_itm;
  wire [286:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  wire [48:0] lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_itm;
  wire [286:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  wire [31:0] lut_lookup_1_else_else_else_else_le_data_f_lshift_1_itm;
  wire [31:0] lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_itm;
  wire mux_3_itm;
  wire mux_20_itm;
  wire mux_25_itm;
  wire mux_26_itm;
  wire mux_582_itm;
  wire mux_595_itm;
  wire mux_tmp_1247;
  wire z_out;
  wire mux_tmp_1250;
  wire z_out_1;
  wire mux_tmp_1253;
  wire z_out_2;
  wire mux_tmp_1257;
  wire and_tmp_201;
  wire z_out_3;
  wire [8:0] z_out_4;
  wire [9:0] nl_z_out_4;
  wire [8:0] z_out_5;
  wire [9:0] nl_z_out_5;
  wire [8:0] z_out_6;
  wire [9:0] nl_z_out_6;
  wire [8:0] z_out_7;
  wire [9:0] nl_z_out_7;
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp;
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp;
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1;
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp_1;
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp_2;
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2;
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3;
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp_3;
  wire chn_lut_in_rsci_ld_core_psct_mx0c0;
  wire main_stage_v_1_mx0c1;
  wire IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0;
  wire FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0;
  wire FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0;
  wire FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0;
  wire FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0;
  wire FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0;
  wire FpMantRNE_49U_24U_1_else_carry_sva_mx0w0;
  wire FpMantRNE_49U_24U_2_else_carry_sva_mx0w0;
  wire main_stage_v_4_mx0c1;
  wire lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1;
  wire lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0;
  wire lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1;
  wire lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0;
  wire lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1;
  wire lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0;
  wire main_stage_v_5_mx0c1;
  wire lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1;
  wire lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1;
  wire lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1;
  wire lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1;
  wire lut_lookup_if_unequal_tmp_1_mx0w0;
  wire lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  wire lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  wire lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  wire lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  wire lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  wire IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0;
  wire [31:0] lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0;
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0;
  wire [31:0] lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0;
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0;
  wire [31:0] lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0;
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0;
  wire [31:0] lut_lookup_if_else_else_le_data_sub_sva_mx0w0;
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_sva_mx0w0;
  wire lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3;
  wire lut_lookup_unequal_tmp_mx0w0;
  wire lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3;
  wire lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3;
  wire lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3;
  wire [22:0] FpAdd_8U_23U_asn_50_mx0w1;
  wire [8:0] lut_lookup_1_else_else_else_else_acc_itm_mx0w0;
  wire [9:0] nl_lut_lookup_1_else_else_else_else_acc_itm_mx0w0;
  wire [22:0] FpAdd_8U_23U_2_asn_50_mx0w1;
  wire [22:0] FpAdd_8U_23U_2_asn_45_mx0w1;
  wire [22:0] FpAdd_8U_23U_2_asn_40_mx0w1;
  wire [22:0] FpAdd_8U_23U_2_asn_35_mx0w1;
  wire IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  wire [22:0] FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_and_tmp;
  wire [22:0] FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_and_tmp;
  wire [22:0] FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_and_1_tmp;
  wire [22:0] FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_and_2_tmp;
  wire [22:0] FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_2_and_3_tmp;
  wire lut_lookup_else_2_else_if_mux_2_cse_mx0;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse;
  wire [34:0] lut_lookup_le_fraction_1_lpi_1_dfm_9;
  wire [8:0] lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1;
  wire [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1;
  wire [34:0] lut_lookup_lo_fraction_1_lpi_1_dfm_1;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse;
  wire lut_lookup_else_2_else_if_mux_7_cse_mx0;
  wire [34:0] lut_lookup_le_fraction_2_lpi_1_dfm_9;
  wire [8:0] lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1;
  wire [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1;
  wire [34:0] lut_lookup_lo_fraction_2_lpi_1_dfm_1;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse;
  wire lut_lookup_else_2_else_if_mux_12_cse_mx0;
  wire [34:0] lut_lookup_le_fraction_3_lpi_1_dfm_9;
  wire [8:0] lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1;
  wire [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1;
  wire [34:0] lut_lookup_lo_fraction_3_lpi_1_dfm_1;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse;
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse;
  wire lut_lookup_else_2_else_if_mux_17_cse_mx0;
  wire [34:0] lut_lookup_le_fraction_lpi_1_dfm_9;
  wire [8:0] lut_lookup_if_1_else_lo_int_lpi_1_dfm_1;
  wire [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_1;
  wire [34:0] lut_lookup_lo_fraction_lpi_1_dfm_1;
  wire lut_lookup_lut_lookup_nor_19_cse;
  wire lut_lookup_and_5_cse;
  wire lut_lookup_and_6_cse;
  wire lut_lookup_and_7_cse;
  wire lut_lookup_lut_lookup_nor_18_cse;
  wire lut_lookup_and_13_cse;
  wire lut_lookup_and_14_cse;
  wire lut_lookup_and_15_cse;
  wire lut_lookup_lut_lookup_nor_17_cse;
  wire lut_lookup_and_21_cse;
  wire lut_lookup_and_22_cse;
  wire lut_lookup_and_23_cse;
  wire lut_lookup_lut_lookup_nor_16_cse;
  wire lut_lookup_and_29_cse;
  wire lut_lookup_and_30_cse;
  wire lut_lookup_and_31_cse;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_1_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_1_sva;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_1_sva;
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_2_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_2_sva;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_2_sva;
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_3_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_3_sva;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_3_sva;
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_sva;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1;
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_sva;
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0;
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva;
  wire [48:0] FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0;
  wire [48:0] FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0;
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva;
  wire [48:0] FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0;
  wire [48:0] FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0;
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva;
  wire [48:0] FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0;
  wire [48:0] FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0;
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva;
  wire [48:0] FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0;
  wire [31:0] lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  wire [32:0] nl_lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  wire [31:0] lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  wire [32:0] nl_lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  wire FpNormalize_8U_49U_oelse_not_9;
  wire FpNormalize_8U_49U_2_oelse_not_9;
  wire FpNormalize_8U_49U_oelse_not_11;
  wire FpNormalize_8U_49U_2_oelse_not_11;
  wire FpNormalize_8U_49U_oelse_not_13;
  wire FpNormalize_8U_49U_2_oelse_not_13;
  wire FpNormalize_8U_49U_oelse_not_15;
  wire FpNormalize_8U_49U_2_oelse_not_15;
  wire [1:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6;
  wire [1:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6;
  wire [1:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6;
  wire [1:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6;
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_4;
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_5;
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_6;
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_7;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19;
  wire [7:0] lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt;
  wire [9:0] nl_lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt;
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire FpAdd_8U_23U_o_expo_and_ssc;
  wire FpAdd_8U_23U_and_57_ssc;
  wire FpAdd_8U_23U_and_49_ssc;
  wire [7:0] lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt;
  wire [9:0] nl_lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt;
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire FpAdd_8U_23U_o_expo_and_1_ssc;
  wire FpAdd_8U_23U_and_55_ssc;
  wire FpAdd_8U_23U_and_47_ssc;
  wire [7:0] lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt;
  wire [9:0] nl_lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt;
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire FpAdd_8U_23U_o_expo_and_2_ssc;
  wire FpAdd_8U_23U_and_53_ssc;
  wire FpAdd_8U_23U_and_45_ssc;
  wire [7:0] lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt;
  wire [9:0] nl_lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt;
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt;
  wire FpAdd_8U_23U_o_expo_and_3_ssc;
  wire FpAdd_8U_23U_and_51_ssc;
  wire FpAdd_8U_23U_and_43_ssc;
  wire cfg_precision_and_cse;
  wire cfg_lut_le_index_offset_and_1_cse;
  wire or_cse;
  wire FpAdd_8U_23U_2_and_35_cse;
  wire FpAdd_8U_23U_2_and_36_cse;
  wire nor_874_cse;
  wire FpAdd_8U_23U_2_and_37_cse;
  wire cfg_lut_le_start_and_cse;
  wire FpMantRNE_49U_24U_1_else_o_mant_and_cse;
  wire nor_5_cse_1;
  wire IsNaN_8U_23U_3_aelse_and_6_cse;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse;
  reg reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  wire FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse;
  wire FpMantRNE_49U_24U_1_else_o_mant_and_1_cse;
  wire nor_27_cse_1;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse;
  reg reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  wire IsNaN_8U_23U_8_aelse_and_1_cse;
  wire FpMantRNE_49U_24U_1_else_o_mant_and_2_cse;
  wire nor_38_cse_1;
  reg reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  wire FpMantRNE_49U_24U_1_else_o_mant_and_3_cse;
  wire nor_50_cse_1;
  reg reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse;
  wire cfg_precision_and_24_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse;
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse;
  wire cfg_lut_hybrid_priority_and_cse;
  wire lut_lookup_lo_index_0_and_cse;
  wire lut_lookup_le_uflow_and_cse;
  wire lut_lookup_else_else_lut_lookup_else_else_or_3_cse;
  wire lut_lookup_lo_index_0_and_2_cse;
  wire lut_lookup_lo_uflow_and_4_cse;
  wire FpAdd_8U_23U_2_is_addition_and_cse;
  wire FpAdd_8U_23U_1_is_addition_and_1_cse;
  reg reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  wire IsZero_8U_23U_4_and_cse;
  wire lut_lookup_FpAdd_8U_23U_1_or_11_cse;
  wire IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse;
  wire lut_lookup_FpAdd_8U_23U_2_or_10_cse;
  wire lut_lookup_FpAdd_8U_23U_2_or_9_cse;
  wire IsZero_8U_23U_7_and_3_cse;
  wire lut_lookup_FpAdd_8U_23U_2_or_8_cse;
  wire IsNaN_8U_23U_3_aelse_and_3_cse;
  wire nor_792_cse;
  wire lut_lookup_lo_index_0_and_4_cse;
  wire lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse;
  wire lut_lookup_lo_index_0_and_6_cse;
  wire lut_lookup_lo_index_0_and_8_cse;
  wire IsNaN_8U_23U_8_and_cse;
  wire IsNaN_8U_23U_8_and_2_cse;
  wire IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse;
  wire and_1142_cse;
  wire nor_832_cse;
  wire and_1138_cse;
  wire and_1139_cse;
  wire and_1140_cse;
  wire and_1141_cse;
  wire or_48_cse;
  wire nor_813_cse;
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse;
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse;
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse;
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse;
  reg [1:0] reg_cfg_precision_1_sva_st_12_cse_1;
  reg reg_cfg_lut_le_function_1_sva_st_19_cse;
  wire and_956_cse;
  wire and_961_cse;
  wire nor_855_cse;
  reg reg_lut_lookup_if_unequal_cse;
  reg reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  reg reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  reg reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  reg reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  reg reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  reg reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  reg reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  wire IsZero_8U_23U_4_and_1_cse;
  wire FpAdd_8U_23U_2_and_44_cse;
  wire lut_lookup_else_and_8_cse;
  wire or_1936_cse;
  reg [1:0] reg_cfg_precision_1_sva_st_13_cse_1;
  reg reg_cfg_lut_le_function_1_sva_st_20_cse;
  wire nor_865_cse;
  wire FpAdd_8U_23U_1_is_a_greater_oelse_and_cse;
  wire FpAdd_8U_23U_2_is_a_greater_oelse_and_cse;
  wire or_849_cse;
  wire nor_190_cse;
  wire mux_580_cse;
  wire or_1688_cse;
  wire nand_95_cse;
  wire nor_196_cse;
  wire mux_1122_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse;
  wire and_401_cse;
  wire FpAdd_8U_23U_1_and_46_cse;
  wire IsNaN_8U_23U_1_aelse_and_5_cse;
  wire IsNaN_8U_23U_1_aelse_and_4_cse;
  wire or_1691_cse;
  wire mux_982_cse;
  wire and_42_cse;
  wire and_832_cse;
  wire nor_193_cse;
  reg reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  wire IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse;
  wire mux_1126_cse;
  wire and_427_cse;
  wire or_312_cse;
  wire IsNaN_8U_23U_7_aelse_and_17_cse;
  wire mux_670_cse;
  wire and_636_cse;
  wire mux_745_cse;
  wire mux_771_cse;
  wire and_898_cse;
  wire and_901_cse;
  wire and_907_cse;
  wire lut_lookup_else_1_and_16_cse;
  wire and_826_cse;
  reg reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  wire FpMantRNE_49U_24U_1_else_and_cse;
  wire mux_83_cse;
  wire lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse;
  wire lut_lookup_if_else_if_and_cse;
  wire FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse;
  wire and_852_cse;
  wire or_492_cse;
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse;
  wire nor_634_cse;
  wire mux_1285_cse;
  wire lut_lookup_if_if_oelse_1_and_cse;
  wire lut_lookup_if_else_if_and_4_cse;
  wire mux_1187_cse;
  wire mux_1188_cse;
  wire and_134_cse;
  wire lut_lookup_else_1_and_13_cse;
  wire FpAdd_8U_23U_2_is_inf_and_cse;
  wire FpAdd_8U_23U_1_is_inf_and_1_cse;
  wire lut_lookup_else_else_and_cse;
  wire lut_lookup_if_1_oelse_1_and_12_cse;
  wire lut_lookup_else_else_and_5_cse;
  wire and_178_cse;
  wire lut_lookup_else_else_and_9_cse;
  wire lut_lookup_else_1_and_9_cse;
  wire and_843_cse;
  wire or_1851_cse;
  wire mux_793_cse;
  wire lut_lookup_if_1_oelse_1_and_4_cse;
  wire lut_lookup_if_1_oelse_1_and_5_cse;
  wire lut_lookup_else_if_oelse_1_and_8_cse;
  wire lut_lookup_if_1_oelse_1_and_14_cse;
  wire mux_805_cse;
  wire lut_lookup_else_1_and_6_cse;
  wire mux_283_cse;
  wire lut_lookup_if_1_oelse_1_and_8_cse;
  wire lut_lookup_else_if_oelse_1_and_1_cse;
  wire lut_lookup_else_if_oelse_1_and_4_cse;
  wire lut_lookup_1_if_else_else_acc_itm_10;
  wire lut_lookup_1_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_2_if_else_else_acc_itm_10;
  wire lut_lookup_2_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_3_if_else_else_acc_itm_10;
  wire lut_lookup_3_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_4_if_else_else_acc_itm_10;
  wire lut_lookup_4_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_1_if_else_else_else_else_acc_itm_32_1;
  wire lut_lookup_1_if_else_else_else_if_acc_itm_3;
  wire lut_lookup_2_if_else_else_else_else_acc_itm_32_1;
  wire lut_lookup_2_if_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_3_if_else_else_else_else_acc_itm_32_1;
  wire lut_lookup_3_if_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_4_if_else_else_else_else_acc_itm_32_1;
  wire lut_lookup_4_if_else_else_else_if_acc_itm_3_1;
  wire lut_lookup_1_else_1_acc_itm_32;
  wire lut_lookup_2_else_1_acc_itm_32;
  wire lut_lookup_3_else_1_acc_itm_32;
  wire lut_lookup_4_else_1_acc_itm_32;
  wire FpAdd_8U_23U_2_is_a_greater_acc_itm_8_1;
  wire FpAdd_8U_23U_2_is_a_greater_acc_1_itm_8_1;
  wire FpAdd_8U_23U_2_is_a_greater_acc_2_itm_8_1;
  wire FpAdd_8U_23U_2_is_a_greater_acc_3_itm_8_1;
  wire lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  wire lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  wire lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  wire lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  wire lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  wire lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  wire lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  wire lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  wire lut_lookup_1_if_if_else_acc_itm_9_1;
  wire lut_lookup_2_if_if_else_acc_itm_9_1;
  wire lut_lookup_3_if_if_else_acc_itm_9_1;
  wire lut_lookup_4_if_if_else_acc_itm_9_1;
  wire lut_lookup_1_else_if_else_if_acc_itm_3_1;
  wire lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  wire lut_lookup_2_else_if_else_if_acc_itm_3_1;
  wire lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  wire lut_lookup_3_else_if_else_if_acc_itm_3_1;
  wire lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  wire lut_lookup_4_else_if_else_if_acc_itm_3_1;
  wire lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  wire lut_lookup_1_if_if_else_else_if_acc_itm_3;
  wire lut_lookup_2_if_if_else_else_if_acc_itm_3;
  wire lut_lookup_3_if_if_else_else_if_acc_itm_3;
  wire lut_lookup_4_if_if_else_else_if_acc_itm_3;
  wire lut_lookup_1_else_else_acc_1_itm_32;
  wire lut_lookup_3_else_else_acc_1_itm_32;
  wire lut_lookup_2_else_else_acc_1_itm_32;
  wire lut_lookup_4_else_else_acc_1_itm_32;
  wire FpAdd_8U_23U_1_is_a_greater_acc_4_itm_8_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_6_itm_8_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_8_itm_8_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_10_itm_8_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1;
  wire lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  wire lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  wire lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  wire lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  wire lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  wire lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  wire lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  wire lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_itm_23_1;
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_itm_23_1;
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_itm_23_1;
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_itm_23_1;
  wire nor_690_cse;
  wire or_365_cse;
  wire mux_851_cse;

  wire[11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_7_nl;
  wire[0:0] lut_lookup_not_39_nl;
  wire[11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_6_nl;
  wire[0:0] lut_lookup_not_38_nl;
  wire[11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_5_nl;
  wire[0:0] lut_lookup_not_37_nl;
  wire[11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_4_nl;
  wire[0:0] lut_lookup_not_36_nl;
  wire[0:0] lut_lookup_else_2_mux_1_nl;
  wire[0:0] lut_lookup_else_2_if_mux_5_nl;
  wire[0:0] lut_lookup_else_2_else_lut_lookup_else_2_else_and_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_61_nl;
  wire[0:0] lut_lookup_else_2_mux_27_nl;
  wire[0:0] lut_lookup_else_2_if_mux_11_nl;
  wire[0:0] lut_lookup_else_2_else_lut_lookup_else_2_else_and_2_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_60_nl;
  wire[0:0] lut_lookup_else_2_mux_53_nl;
  wire[0:0] lut_lookup_else_2_if_mux_17_nl;
  wire[0:0] lut_lookup_else_2_else_lut_lookup_else_2_else_and_4_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_59_nl;
  wire[0:0] lut_lookup_else_2_mux_79_nl;
  wire[0:0] lut_lookup_else_2_if_mux_23_nl;
  wire[0:0] lut_lookup_else_2_else_lut_lookup_else_2_else_and_6_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_nl;
  wire[0:0] lut_lookup_else_2_lut_lookup_else_2_and_4_nl;
  wire[0:0] lut_lookup_else_2_lut_lookup_else_2_and_5_nl;
  wire[0:0] lut_lookup_else_2_lut_lookup_else_2_and_6_nl;
  wire[0:0] lut_lookup_else_2_lut_lookup_else_2_and_7_nl;
  wire[0:0] lut_lookup_else_2_mux_103_nl;
  wire[0:0] lut_lookup_else_2_else_mux_3_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_3_nl;
  wire[0:0] lut_lookup_else_2_mux_104_nl;
  wire[0:0] lut_lookup_else_2_else_mux_23_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_18_nl;
  wire[0:0] lut_lookup_else_2_mux_105_nl;
  wire[0:0] lut_lookup_else_2_else_mux_43_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_33_nl;
  wire[0:0] lut_lookup_else_2_mux_106_nl;
  wire[0:0] lut_lookup_else_2_else_mux_63_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_48_nl;
  wire[5:0] lut_lookup_else_if_lut_lookup_else_if_and_2_nl;
  wire[0:0] lut_lookup_else_2_mux_107_nl;
  wire[0:0] lut_lookup_else_2_else_mux_18_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_13_nl;
  wire[0:0] lut_lookup_if_2_mux_21_nl;
  wire[0:0] lut_lookup_else_2_mux_108_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_1_nl;
  wire[0:0] lut_lookup_else_2_else_mux_17_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_12_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_3_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_8_nl;
  wire[0:0] lut_lookup_else_2_mux_109_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_nl;
  wire[0:0] lut_lookup_else_2_else_mux_16_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_11_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_2_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_9_nl;
  wire[5:0] lut_lookup_else_if_lut_lookup_else_if_and_5_nl;
  wire[0:0] lut_lookup_else_2_mux_110_nl;
  wire[0:0] lut_lookup_else_2_else_mux_38_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_28_nl;
  wire[0:0] lut_lookup_if_2_mux_22_nl;
  wire[0:0] lut_lookup_else_2_mux_111_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_3_nl;
  wire[0:0] lut_lookup_else_2_else_mux_37_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_27_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_7_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_10_nl;
  wire[0:0] lut_lookup_else_2_mux_112_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_2_nl;
  wire[0:0] lut_lookup_else_2_else_mux_36_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_26_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_6_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_11_nl;
  wire[5:0] lut_lookup_else_if_lut_lookup_else_if_and_8_nl;
  wire[0:0] lut_lookup_else_2_mux_113_nl;
  wire[0:0] lut_lookup_else_2_else_mux_58_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_43_nl;
  wire[0:0] lut_lookup_if_2_mux_23_nl;
  wire[0:0] lut_lookup_else_2_mux_114_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_5_nl;
  wire[0:0] lut_lookup_else_2_else_mux_57_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_42_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_11_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_12_nl;
  wire[0:0] lut_lookup_else_2_mux_115_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_4_nl;
  wire[0:0] lut_lookup_else_2_else_mux_56_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_41_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_10_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_13_nl;
  wire[5:0] lut_lookup_else_if_lut_lookup_else_if_and_11_nl;
  wire[0:0] lut_lookup_else_2_mux_116_nl;
  wire[0:0] lut_lookup_else_2_else_mux_78_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_58_nl;
  wire[0:0] lut_lookup_if_2_mux_24_nl;
  wire[0:0] lut_lookup_else_2_mux_117_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_7_nl;
  wire[0:0] lut_lookup_else_2_else_mux_77_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_57_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_15_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_14_nl;
  wire[0:0] lut_lookup_else_2_mux_118_nl;
  wire[0:0] lut_lookup_else_2_if_lut_lookup_else_2_if_and_6_nl;
  wire[0:0] lut_lookup_else_2_else_mux_76_nl;
  wire[0:0] lut_lookup_else_2_else_else_mux_56_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_14_nl;
  wire[0:0] lut_lookup_if_2_lut_lookup_if_2_and_15_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] nor_783_nl;
  wire[49:0] lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[49:0] lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl;
  wire[49:0] lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl;
  wire[49:0] lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[49:0] lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[49:0] lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[49:0] lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl;
  wire[49:0] lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl;
  wire[49:0] lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[49:0] lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[49:0] lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[49:0] lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl;
  wire[49:0] lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl;
  wire[49:0] lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[49:0] lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[49:0] lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[49:0] lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl;
  wire[49:0] lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl;
  wire[49:0] lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[50:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl;
  wire[49:0] lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[51:0] nl_lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] or_2081_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] or_1931_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] mux_1220_nl;
  wire[1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl;
  wire[5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl;
  wire[0:0] FpAdd_8U_23U_o_expo_or_3_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] or_1941_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] and_868_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] and_869_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] nor_773_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] and_45_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] nor_770_nl;
  wire[7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_nl;
  wire[7:0] lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl;
  wire[9:0] nl_lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] or_114_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] or_118_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] or_120_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] or_125_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] or_40_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] or_2080_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] or_1948_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] mux_1227_nl;
  wire[1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl;
  wire[5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_10_nl;
  wire[0:0] FpAdd_8U_23U_o_expo_or_2_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] nor_852_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] and_864_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] and_865_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_760_nl;
  wire[0:0] nor_761_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] nor_757_nl;
  wire[0:0] and_48_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] nor_758_nl;
  wire[7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_2_nl;
  wire[7:0] lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl;
  wire[9:0] nl_lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] and_49_nl;
  wire[0:0] or_184_nl;
  wire[0:0] nor_35_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] or_2079_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] or_1964_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] nor_749_nl;
  wire[0:0] nor_750_nl;
  wire[1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl;
  wire[0:0] mux_1233_nl;
  wire[5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl;
  wire[0:0] FpAdd_8U_23U_o_expo_or_1_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] or_1976_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] and_861_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] and_862_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] nor_745_nl;
  wire[0:0] nor_746_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] nor_742_nl;
  wire[0:0] and_54_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] nor_743_nl;
  wire[7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_4_nl;
  wire[7:0] lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl;
  wire[9:0] nl_lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] or_247_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] or_251_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] or_2078_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] or_1983_nl;
  wire[0:0] nor_802_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] nor_737_nl;
  wire[0:0] nor_738_nl;
  wire[1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl;
  wire[0:0] mux_1240_nl;
  wire[5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_8_nl;
  wire[0:0] FpAdd_8U_23U_o_expo_or_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] or_1995_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] and_858_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] and_859_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] and_59_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] nor_730_nl;
  wire[7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_6_nl;
  wire[7:0] lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl;
  wire[9:0] nl_lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] nand_76_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] or_306_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] or_311_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] or_315_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] nor_726_nl;
  wire[0:0] nor_727_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] nor_724_nl;
  wire[0:0] nor_725_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] nor_722_nl;
  wire[0:0] nor_723_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] and_62_nl;
  wire[0:0] nor_721_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] or_332_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_63_nl;
  wire[0:0] and_64_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] or_341_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] or_346_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] nor_719_nl;
  wire[0:0] nor_720_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] nor_715_nl;
  wire[0:0] nor_716_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] nor_713_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] and_69_nl;
  wire[0:0] nor_714_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] and_70_nl;
  wire[0:0] and_71_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] or_374_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] nor_712_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] nor_708_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] and_74_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] and_75_nl;
  wire[0:0] and_76_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] or_406_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] or_411_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] nor_705_nl;
  wire[0:0] nor_706_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] nor_701_nl;
  wire[0:0] nor_702_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] and_79_nl;
  wire[0:0] nor_700_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] and_80_nl;
  wire[0:0] and_81_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] and_447_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] nor_698_nl;
  wire[0:0] nor_699_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] nor_697_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] or_445_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] or_475_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] and_451_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] or_528_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] and_455_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] or_545_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] or_566_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] or_569_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] or_575_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] and_459_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] or_596_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] or_617_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] or_620_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] or_625_nl;
  wire[34:0] lut_lookup_if_else_else_else_else_mux_nl;
  wire[34:0] lut_lookup_if_else_else_else_else_mux_1_nl;
  wire[34:0] lut_lookup_if_else_else_else_else_mux_2_nl;
  wire[34:0] lut_lookup_if_else_else_else_else_mux_3_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] lut_lookup_else_else_lut_lookup_else_else_and_10_nl;
  wire[0:0] lut_lookup_if_else_lut_lookup_if_else_and_11_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_4_nl;
  wire[0:0] lut_lookup_else_else_lut_lookup_else_else_and_7_nl;
  wire[0:0] lut_lookup_if_else_lut_lookup_if_else_and_12_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_5_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] lut_lookup_else_else_lut_lookup_else_else_and_4_nl;
  wire[0:0] lut_lookup_if_else_lut_lookup_if_else_and_13_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_6_nl;
  wire[0:0] lut_lookup_else_else_lut_lookup_else_else_and_1_nl;
  wire[0:0] lut_lookup_if_else_lut_lookup_if_else_and_14_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_7_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] and_830_nl;
  wire[0:0] mux_371_nl;
  wire[8:0] acc_4_nl;
  wire[9:0] nl_acc_4_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_8_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_9_nl;
  wire[8:0] acc_6_nl;
  wire[9:0] nl_acc_6_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_10_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_11_nl;
  wire[8:0] acc_8_nl;
  wire[9:0] nl_acc_8_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_12_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_13_nl;
  wire[8:0] acc_10_nl;
  wire[9:0] nl_acc_10_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_14_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_15_nl;
  wire[8:0] acc_11_nl;
  wire[9:0] nl_acc_11_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_14_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_15_nl;
  wire[8:0] acc_9_nl;
  wire[9:0] nl_acc_9_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_12_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_13_nl;
  wire[8:0] acc_7_nl;
  wire[9:0] nl_acc_7_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_10_nl;
  wire[7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_11_nl;
  wire[8:0] acc_5_nl;
  wire[9:0] nl_acc_5_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_8_nl;
  wire[7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_9_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] or_827_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] or_829_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] or_839_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] or_850_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] or_1696_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] nand_16_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] and_827_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] and_98_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_655_nl;
  wire[0:0] and_100_nl;
  wire[0:0] and_101_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] and_102_nl;
  wire[0:0] and_103_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] and_104_nl;
  wire[0:0] and_105_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] and_106_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] and_108_nl;
  wire[0:0] and_109_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] and_110_nl;
  wire[0:0] and_111_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] and_112_nl;
  wire[0:0] mux_663_nl;
  wire[0:0] or_879_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] or_880_nl;
  wire[0:0] and_113_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] or_885_nl;
  wire[0:0] or_887_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] or_888_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] and_114_nl;
  wire[0:0] mux_674_nl;
  wire[0:0] or_899_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] or_900_nl;
  wire[0:0] and_115_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] mux_675_nl;
  wire[0:0] nand_18_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] or_907_nl;
  wire[0:0] mux_689_nl;
  wire[0:0] and_116_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] or_915_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] or_916_nl;
  wire[0:0] and_117_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] mux_686_nl;
  wire[0:0] nand_19_nl;
  wire[0:0] mux_687_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] or_923_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] and_118_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] or_931_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] or_932_nl;
  wire[0:0] and_119_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] or_939_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] mux_707_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] and_120_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] and_823_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] mux_722_nl;
  wire[0:0] and_822_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] mux_731_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] mux_743_nl;
  wire[0:0] mux_749_nl;
  wire[0:0] mux_748_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] and_1166_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] or_990_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] and_1164_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] and_127_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] and_819_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] mux_774_nl;
  wire[0:0] mux_773_nl;
  wire[0:0] mux_772_nl;
  wire[0:0] nor_609_nl;
  wire[30:0] lut_lookup_1_IntLog2_32U_and_nl;
  wire[30:0] lut_lookup_1_IntLog2_32U_acc_1_nl;
  wire[31:0] nl_lut_lookup_1_IntLog2_32U_acc_1_nl;
  wire[22:0] lut_lookup_lut_lookup_mux_17_nl;
  wire[0:0] and_649_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] and_815_nl;
  wire[0:0] and_816_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] and_131_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] nor_435_nl;
  wire[6:0] lut_lookup_1_if_else_else_else_else_else_acc_nl;
  wire[7:0] nl_lut_lookup_1_if_else_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_1_if_else_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_1_if_else_else_else_else_if_acc_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] and_132_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] or_1045_nl;
  wire[8:0] lut_lookup_1_else_1_else_else_acc_nl;
  wire[9:0] nl_lut_lookup_1_else_1_else_else_acc_nl;
  wire[7:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl;
  wire[8:0] nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] or_2009_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] nor_830_nl;
  wire[0:0] or_2007_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] and_1162_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] or_1072_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] and_1160_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] and_138_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] and_812_nl;
  wire[30:0] lut_lookup_2_IntLog2_32U_and_nl;
  wire[30:0] lut_lookup_2_IntLog2_32U_acc_1_nl;
  wire[31:0] nl_lut_lookup_2_IntLog2_32U_acc_1_nl;
  wire[22:0] lut_lookup_lut_lookup_mux_nl;
  wire[0:0] and_657_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] and_142_nl;
  wire[6:0] lut_lookup_2_if_else_else_else_else_else_acc_nl;
  wire[7:0] nl_lut_lookup_2_if_else_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_2_if_else_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_2_if_else_else_else_else_if_acc_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] and_143_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] or_1113_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] and_1089_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] and_147_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] or_1142_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] and_1156_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] and_149_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] and_808_nl;
  wire[30:0] lut_lookup_3_IntLog2_32U_and_nl;
  wire[30:0] lut_lookup_3_IntLog2_32U_acc_1_nl;
  wire[31:0] nl_lut_lookup_3_IntLog2_32U_acc_1_nl;
  wire[22:0] lut_lookup_lut_lookup_mux_3_nl;
  wire[0:0] and_665_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] and_152_nl;
  wire[6:0] lut_lookup_3_if_else_else_else_else_else_acc_nl;
  wire[7:0] nl_lut_lookup_3_if_else_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_3_if_else_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_3_if_else_else_else_else_if_acc_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] and_153_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] or_1183_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] nor_827_nl;
  wire[0:0] nand_102_nl;
  wire[0:0] or_2025_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] and_158_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] and_1176_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] nor_544_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] and_1153_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] or_1213_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] and_1151_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] and_160_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] and_804_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] and_1174_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] or_2087_nl;
  wire[30:0] lut_lookup_4_IntLog2_32U_and_nl;
  wire[30:0] lut_lookup_4_IntLog2_32U_acc_1_nl;
  wire[31:0] nl_lut_lookup_4_IntLog2_32U_acc_1_nl;
  wire[22:0] lut_lookup_lut_lookup_mux_4_nl;
  wire[0:0] and_672_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] and_163_nl;
  wire[6:0] lut_lookup_4_if_else_else_else_else_else_acc_nl;
  wire[7:0] nl_lut_lookup_4_if_else_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_4_if_else_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_4_if_else_else_else_else_if_acc_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] and_164_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] and_166_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] or_1252_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] nand_nl;
  wire[0:0] or_2035_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] nor_315_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] and_1147_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] and_179_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] and_1179_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] and_1149_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] and_193_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] and_1148_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] and_204_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] and_1146_nl;
  wire[0:0] mux_nl;
  wire[0:0] and_215_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] mux_1061_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_1_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] and_219_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] and_220_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] and_221_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] or_1431_nl;
  wire[5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_3_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] and_222_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] and_224_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] and_226_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] or_1440_nl;
  wire[5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_5_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] and_228_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] and_230_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] and_232_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] or_1450_nl;
  wire[5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_7_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] and_233_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] and_235_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] and_236_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] or_1458_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] or_1460_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] and_774_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] and_773_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] mux_1118_nl;
  wire[10:0] lut_lookup_1_if_else_else_acc_nl;
  wire[11:0] nl_lut_lookup_1_if_else_else_acc_nl;
  wire[3:0] lut_lookup_1_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_1_else_else_else_if_acc_nl;
  wire[10:0] lut_lookup_2_if_else_else_acc_nl;
  wire[11:0] nl_lut_lookup_2_if_else_else_acc_nl;
  wire[3:0] lut_lookup_2_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_2_else_else_else_if_acc_nl;
  wire[10:0] lut_lookup_3_if_else_else_acc_nl;
  wire[11:0] nl_lut_lookup_3_if_else_else_acc_nl;
  wire[3:0] lut_lookup_3_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_3_else_else_else_if_acc_nl;
  wire[10:0] lut_lookup_4_if_else_else_acc_nl;
  wire[11:0] nl_lut_lookup_4_if_else_else_acc_nl;
  wire[3:0] lut_lookup_4_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_4_else_else_else_if_acc_nl;
  wire[32:0] lut_lookup_1_if_else_else_else_else_acc_nl;
  wire[33:0] nl_lut_lookup_1_if_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_1_if_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_1_if_else_else_else_if_acc_nl;
  wire[32:0] lut_lookup_2_if_else_else_else_else_acc_nl;
  wire[33:0] nl_lut_lookup_2_if_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_2_if_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_2_if_else_else_else_if_acc_nl;
  wire[32:0] lut_lookup_3_if_else_else_else_else_acc_nl;
  wire[33:0] nl_lut_lookup_3_if_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_3_if_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_3_if_else_else_else_if_acc_nl;
  wire[32:0] lut_lookup_4_if_else_else_else_else_acc_nl;
  wire[33:0] nl_lut_lookup_4_if_else_else_else_else_acc_nl;
  wire[3:0] lut_lookup_4_if_else_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_4_if_else_else_else_if_acc_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_or_3_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_or_2_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_or_1_nl;
  wire[0:0] lut_lookup_if_if_lut_lookup_if_if_or_nl;
  wire[32:0] lut_lookup_1_else_1_acc_nl;
  wire[33:0] nl_lut_lookup_1_else_1_acc_nl;
  wire[32:0] lut_lookup_2_else_1_acc_nl;
  wire[33:0] nl_lut_lookup_2_else_1_acc_nl;
  wire[32:0] lut_lookup_3_else_1_acc_nl;
  wire[33:0] nl_lut_lookup_3_else_1_acc_nl;
  wire[32:0] lut_lookup_4_else_1_acc_nl;
  wire[33:0] nl_lut_lookup_4_else_1_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl;
  wire[22:0] lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_4_nl;
  wire[22:0] lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[23:0] nl_lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl;
  wire[22:0] lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_5_nl;
  wire[22:0] lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[23:0] nl_lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl;
  wire[22:0] lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_6_nl;
  wire[22:0] lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[23:0] nl_lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl;
  wire[22:0] lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_7_nl;
  wire[22:0] lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[23:0] nl_lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl;
  wire[8:0] FpAdd_8U_23U_2_is_a_greater_acc_nl;
  wire[10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_nl;
  wire[8:0] FpAdd_8U_23U_2_is_a_greater_acc_1_nl;
  wire[10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_2_is_a_greater_acc_2_nl;
  wire[10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_2_nl;
  wire[8:0] FpAdd_8U_23U_2_is_a_greater_acc_3_nl;
  wire[10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_3_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_59_nl;
  wire[0:0] FpAdd_8U_23U_and_61_nl;
  wire[0:0] FpAdd_8U_23U_1_and_35_nl;
  wire[0:0] FpAdd_8U_23U_and_35_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_4_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_2_and_nl;
  wire[0:0] FpAdd_8U_23U_2_and_6_nl;
  wire[0:0] FpAdd_8U_23U_2_and_28_nl;
  wire[0:0] FpAdd_8U_23U_2_and_9_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_63_nl;
  wire[0:0] FpAdd_8U_23U_and_65_nl;
  wire[0:0] FpAdd_8U_23U_1_and_37_nl;
  wire[0:0] FpAdd_8U_23U_and_37_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_5_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_2_and_29_nl;
  wire[0:0] FpAdd_8U_23U_2_and_13_nl;
  wire[0:0] FpAdd_8U_23U_2_and_30_nl;
  wire[0:0] FpAdd_8U_23U_2_and_15_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_67_nl;
  wire[0:0] FpAdd_8U_23U_and_69_nl;
  wire[0:0] FpAdd_8U_23U_1_and_39_nl;
  wire[0:0] FpAdd_8U_23U_and_39_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_6_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_2_and_31_nl;
  wire[0:0] FpAdd_8U_23U_2_and_19_nl;
  wire[0:0] FpAdd_8U_23U_2_and_32_nl;
  wire[0:0] FpAdd_8U_23U_2_and_21_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_71_nl;
  wire[0:0] FpAdd_8U_23U_and_73_nl;
  wire[0:0] FpAdd_8U_23U_1_and_41_nl;
  wire[0:0] FpAdd_8U_23U_and_41_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_7_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_2_and_33_nl;
  wire[0:0] FpAdd_8U_23U_2_and_25_nl;
  wire[0:0] FpAdd_8U_23U_2_and_34_nl;
  wire[0:0] FpAdd_8U_23U_2_and_27_nl;
  wire[9:0] lut_lookup_1_if_if_else_acc_nl;
  wire[10:0] nl_lut_lookup_1_if_if_else_acc_nl;
  wire[9:0] lut_lookup_2_if_if_else_acc_nl;
  wire[10:0] nl_lut_lookup_2_if_if_else_acc_nl;
  wire[9:0] lut_lookup_3_if_if_else_acc_nl;
  wire[10:0] nl_lut_lookup_3_if_if_else_acc_nl;
  wire[9:0] lut_lookup_4_if_if_else_acc_nl;
  wire[10:0] nl_lut_lookup_4_if_if_else_acc_nl;
  wire[3:0] lut_lookup_1_else_if_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_1_else_if_else_if_acc_nl;
  wire[0:0] lut_lookup_else_mux_172_nl;
  wire[0:0] lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_nl;
  wire[0:0] lut_lookup_if_1_lut_lookup_if_1_and_11_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_nl;
  wire[247:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[247:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_nl;
  wire[3:0] lut_lookup_2_else_if_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_2_else_if_else_if_acc_nl;
  wire[0:0] lut_lookup_else_mux_174_nl;
  wire[0:0] lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_1_nl;
  wire[0:0] lut_lookup_if_1_lut_lookup_if_1_and_12_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_1_nl;
  wire[247:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[247:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_1_nl;
  wire[3:0] lut_lookup_3_else_if_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_3_else_if_else_if_acc_nl;
  wire[0:0] lut_lookup_else_mux_176_nl;
  wire[0:0] lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_2_nl;
  wire[0:0] lut_lookup_if_1_lut_lookup_if_1_and_13_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_2_nl;
  wire[247:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[247:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_2_nl;
  wire[3:0] lut_lookup_4_else_if_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_4_else_if_else_if_acc_nl;
  wire[0:0] lut_lookup_if_1_lut_lookup_if_1_and_14_nl;
  wire[0:0] lut_lookup_else_mux_178_nl;
  wire[0:0] lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_3_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_3_nl;
  wire[247:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  wire[247:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[248:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  wire[8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_3_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_30_nl;
  wire[0:0] FpAdd_8U_23U_2_is_a_greater_oelse_not_23_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_32_nl;
  wire[0:0] FpAdd_8U_23U_2_is_a_greater_oelse_not_25_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_34_nl;
  wire[0:0] FpAdd_8U_23U_2_is_a_greater_oelse_not_27_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_36_nl;
  wire[0:0] FpAdd_8U_23U_2_is_a_greater_oelse_not_29_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  wire[0:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_1_nl;
  wire[0:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  wire[0:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_3_nl;
  wire[0:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  wire[0:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_5_nl;
  wire[0:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  wire[0:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  wire[48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_7_nl;
  wire[0:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  wire[3:0] lut_lookup_1_if_if_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_1_if_if_else_else_if_acc_nl;
  wire[3:0] lut_lookup_2_if_if_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_2_if_if_else_else_if_acc_nl;
  wire[3:0] lut_lookup_3_if_if_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_3_if_if_else_else_if_acc_nl;
  wire[3:0] lut_lookup_4_if_if_else_else_if_acc_nl;
  wire[4:0] nl_lut_lookup_4_if_if_else_else_if_acc_nl;
  wire[32:0] lut_lookup_1_else_else_acc_1_nl;
  wire[33:0] nl_lut_lookup_1_else_else_acc_1_nl;
  wire[32:0] lut_lookup_3_else_else_acc_1_nl;
  wire[33:0] nl_lut_lookup_3_else_else_acc_1_nl;
  wire[32:0] lut_lookup_2_else_else_acc_1_nl;
  wire[33:0] nl_lut_lookup_2_else_else_acc_1_nl;
  wire[32:0] lut_lookup_4_else_else_acc_1_nl;
  wire[33:0] nl_lut_lookup_4_else_else_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_4_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_4_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_6_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_6_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_8_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_8_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_10_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_10_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  wire[8:0] lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl;
  wire[10:0] nl_lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl;
  wire[8:0] lut_lookup_1_FpNormalize_8U_49U_2_acc_nl;
  wire[10:0] nl_lut_lookup_1_FpNormalize_8U_49U_2_acc_nl;
  wire[8:0] lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl;
  wire[10:0] nl_lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl;
  wire[8:0] lut_lookup_2_FpNormalize_8U_49U_2_acc_nl;
  wire[10:0] nl_lut_lookup_2_FpNormalize_8U_49U_2_acc_nl;
  wire[8:0] lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl;
  wire[10:0] nl_lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl;
  wire[8:0] lut_lookup_3_FpNormalize_8U_49U_2_acc_nl;
  wire[10:0] nl_lut_lookup_3_FpNormalize_8U_49U_2_acc_nl;
  wire[8:0] lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl;
  wire[10:0] nl_lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl;
  wire[8:0] lut_lookup_4_FpNormalize_8U_49U_2_acc_nl;
  wire[10:0] nl_lut_lookup_4_FpNormalize_8U_49U_2_acc_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  wire[0:0] or_4_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] or_122_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] or_121_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] or_127_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] or_126_nl;
  wire[0:0] nand_93_nl;
  wire[0:0] or_191_nl;
  wire[0:0] or_186_nl;
  wire[0:0] or_302_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] or_1860_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] or_841_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] or_832_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] or_856_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] or_1583_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] or_1594_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] or_1606_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] or_1618_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_1179_nl;
  wire[23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl;
  wire[25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl;
  wire[23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl;
  wire[25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl;
  wire[23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl;
  wire[25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl;
  wire[23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl;
  wire[25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] or_1972_nl;
  wire[0:0] or_1973_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] or_1991_nl;
  wire[0:0] or_1992_nl;
  wire[0:0] nor_823_nl;
  wire[0:0] nor_820_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] or_2056_nl;
  wire[0:0] or_2055_nl;
  wire[0:0] nor_814_nl;
  wire[0:0] lut_lookup_else_2_if_mux_31_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_and_4_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] or_2088_nl;
  wire[0:0] nand_114_nl;
  wire[0:0] lut_lookup_else_2_if_mux_32_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_and_5_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] nand_115_nl;
  wire[0:0] or_2089_nl;
  wire[0:0] nand_116_nl;
  wire[0:0] lut_lookup_else_2_if_mux_33_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_and_6_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] nand_117_nl;
  wire[0:0] or_2090_nl;
  wire[0:0] nand_118_nl;
  wire[0:0] lut_lookup_else_2_if_mux_34_nl;
  wire[0:0] lut_lookup_else_2_else_else_else_and_7_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] nor_882_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm};
  wire [9:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s = (lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm};
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = {1'b1
      , FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5};
  wire [9:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = (lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a =
      {1'b1 , FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5};
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg};
  wire [9:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s = (lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg};
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = {1'b1
      , FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5};
  wire [9:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = (lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a =
      {1'b1 , FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5};
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg};
  wire [9:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s = (lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg};
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = {1'b1
      , FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5};
  wire [9:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = (lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a =
      {1'b1 , FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5};
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1};
  wire [9:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s = (lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = {1'b1
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1};
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = {1'b1
      , FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5};
  wire [9:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = (lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0])
      + 9'b100011;
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a =
      {1'b1 , FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5};
  wire [30:0] nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_a;
  assign nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm};
  wire [5:0] nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_s;
  assign nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_s = {reg_lut_lookup_1_else_else_else_else_acc_3_reg
      , lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3};
  wire [30:0] nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm};
  wire [7:0] nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_s = {1'b1 , reg_lut_lookup_1_else_else_else_else_acc_2_reg
      , reg_lut_lookup_1_else_else_else_else_acc_3_reg};
  wire [34:0] nl_lut_lookup_1_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_1_else_else_else_else_rshift_rg_a = {{3{lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31]}},
      lut_lookup_1_else_else_else_else_le_data_f_and_itm_2};
  wire [8:0] nl_lut_lookup_1_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_1_else_else_else_else_rshift_rg_s = {reg_lut_lookup_1_else_else_else_else_acc_reg
      , reg_lut_lookup_1_else_else_else_else_acc_1_reg , reg_lut_lookup_1_else_else_else_else_acc_2_reg
      , reg_lut_lookup_1_else_else_else_else_acc_3_reg};
  wire [8:0] nl_lut_lookup_1_else_1_else_else_rshift_rg_s;
  assign nl_lut_lookup_1_else_1_else_else_rshift_rg_s = {reg_lut_lookup_1_else_1_else_else_acc_itm
      , reg_lut_lookup_1_else_1_else_else_acc_1_itm};
  wire [30:0] nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_a;
  assign nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg};
  wire [5:0] nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_s;
  assign nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_s = {reg_lut_lookup_2_else_else_else_else_acc_3_reg
      , lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3};
  wire [30:0] nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg};
  wire [7:0] nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_s = {1'b1 , reg_lut_lookup_2_else_else_else_else_acc_2_reg
      , reg_lut_lookup_2_else_else_else_else_acc_3_reg};
  wire [34:0] nl_lut_lookup_2_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_2_else_else_else_else_rshift_rg_a = {{3{lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31]}},
      lut_lookup_2_else_else_else_else_le_data_f_and_itm_2};
  wire [8:0] nl_lut_lookup_2_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_2_else_else_else_else_rshift_rg_s = {reg_lut_lookup_2_else_else_else_else_acc_reg
      , reg_lut_lookup_2_else_else_else_else_acc_1_reg , reg_lut_lookup_2_else_else_else_else_acc_2_reg
      , reg_lut_lookup_2_else_else_else_else_acc_3_reg};
  wire [8:0] nl_lut_lookup_2_else_1_else_else_rshift_rg_s;
  assign nl_lut_lookup_2_else_1_else_else_rshift_rg_s = {reg_lut_lookup_2_else_1_else_else_acc_itm
      , reg_lut_lookup_2_else_1_else_else_acc_1_itm};
  wire [30:0] nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_a;
  assign nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg};
  wire [5:0] nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_s;
  assign nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_s = {reg_lut_lookup_3_else_else_else_else_acc_3_reg
      , lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3};
  wire [30:0] nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg};
  wire [7:0] nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_s = {1'b1 , reg_lut_lookup_3_else_else_else_else_acc_2_reg
      , reg_lut_lookup_3_else_else_else_else_acc_3_reg};
  wire [34:0] nl_lut_lookup_3_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_3_else_else_else_else_rshift_rg_a = {{3{lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31]}},
      lut_lookup_3_else_else_else_else_le_data_f_and_itm_2};
  wire [8:0] nl_lut_lookup_3_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_3_else_else_else_else_rshift_rg_s = {reg_lut_lookup_3_else_else_else_else_acc_reg
      , reg_lut_lookup_3_else_else_else_else_acc_1_reg , reg_lut_lookup_3_else_else_else_else_acc_2_reg
      , reg_lut_lookup_3_else_else_else_else_acc_3_reg};
  wire [8:0] nl_lut_lookup_3_else_1_else_else_rshift_rg_s;
  assign nl_lut_lookup_3_else_1_else_else_rshift_rg_s = {reg_lut_lookup_3_else_1_else_else_acc_itm
      , reg_lut_lookup_3_else_1_else_else_acc_1_itm};
  wire [30:0] nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_a;
  assign nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_reg
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1};
  wire [5:0] nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_s;
  assign nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_s = {reg_lut_lookup_4_else_else_else_else_acc_3_reg
      , lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3};
  wire [30:0] nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_a = {reg_IntLog2_32U_ac_int_cctor_1_30_0_reg
      , reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1};
  wire [7:0] nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_s = {1'b1 , reg_lut_lookup_4_else_else_else_else_acc_2_reg
      , reg_lut_lookup_4_else_else_else_else_acc_3_reg};
  wire [34:0] nl_lut_lookup_4_else_else_else_else_rshift_rg_a;
  assign nl_lut_lookup_4_else_else_else_else_rshift_rg_a = {{3{lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31]}},
      lut_lookup_4_else_else_else_else_le_data_f_and_itm_2};
  wire [8:0] nl_lut_lookup_4_else_else_else_else_rshift_rg_s;
  assign nl_lut_lookup_4_else_else_else_else_rshift_rg_s = {reg_lut_lookup_4_else_else_else_else_acc_reg
      , reg_lut_lookup_4_else_else_else_else_acc_1_reg , reg_lut_lookup_4_else_else_else_else_acc_2_reg
      , reg_lut_lookup_4_else_else_else_else_acc_3_reg};
  wire [8:0] nl_lut_lookup_4_else_1_else_else_rshift_rg_s;
  assign nl_lut_lookup_4_else_1_else_else_rshift_rg_s = {reg_lut_lookup_4_else_1_else_else_acc_itm
      , reg_lut_lookup_4_else_1_else_else_acc_1_itm};
  wire [31:0] nl_lut_lookup_1_IntLog2_32U_lshift_rg_s;
  assign nl_lut_lookup_1_IntLog2_32U_lshift_rg_s = signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[4:0]))});
  wire [31:0] nl_lut_lookup_2_IntLog2_32U_lshift_rg_s;
  assign nl_lut_lookup_2_IntLog2_32U_lshift_rg_s = signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[4:0]))});
  wire [31:0] nl_lut_lookup_3_IntLog2_32U_lshift_rg_s;
  assign nl_lut_lookup_3_IntLog2_32U_lshift_rg_s = signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[4:0]))});
  wire [31:0] nl_lut_lookup_4_IntLog2_32U_lshift_rg_s;
  assign nl_lut_lookup_4_IntLog2_32U_lshift_rg_s = signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[4:0]))});
  wire [48:0] nl_lut_lookup_1_leading_sign_49_0_rg_mantissa;
  assign nl_lut_lookup_1_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  wire [48:0] nl_lut_lookup_1_leading_sign_49_0_2_rg_mantissa;
  assign nl_lut_lookup_1_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0];
  wire [48:0] nl_lut_lookup_2_leading_sign_49_0_rg_mantissa;
  assign nl_lut_lookup_2_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  wire [48:0] nl_lut_lookup_2_leading_sign_49_0_2_rg_mantissa;
  assign nl_lut_lookup_2_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0];
  wire [48:0] nl_lut_lookup_3_leading_sign_49_0_rg_mantissa;
  assign nl_lut_lookup_3_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  wire [48:0] nl_lut_lookup_3_leading_sign_49_0_2_rg_mantissa;
  assign nl_lut_lookup_3_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0];
  wire [48:0] nl_lut_lookup_4_leading_sign_49_0_rg_mantissa;
  assign nl_lut_lookup_4_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  wire [48:0] nl_lut_lookup_4_leading_sign_49_0_2_rg_mantissa;
  assign nl_lut_lookup_4_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0];
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (lut_in_data_sva_154[22:0])};
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (lut_in_data_sva_154[22:0])};
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2
      , (cfg_lut_lo_start_1_sva_41[22:0])};
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s = {(lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = {lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2
      , (lut_in_data_sva_154[22:0])};
  wire[7:0] lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s = {(lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (lut_in_data_sva_154[54:32])};
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (lut_in_data_sva_154[54:32])};
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2
      , (cfg_lut_lo_start_1_sva_41[22:0])};
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s = {(lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = {lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2
      , (lut_in_data_sva_154[54:32])};
  wire[7:0] lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s = {(lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (lut_in_data_sva_154[86:64])};
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (lut_in_data_sva_154[86:64])};
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2
      , (cfg_lut_lo_start_1_sva_41[22:0])};
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s = {(lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = {lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2
      , (lut_in_data_sva_154[86:64])};
  wire[7:0] lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s = {(lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (lut_in_data_sva_154[118:96])};
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2
      , (cfg_lut_le_start_1_sva_41[22:0])};
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , (lut_in_data_sva_154[118:96])};
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1
      , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2
      , (cfg_lut_lo_start_1_sva_41[22:0])};
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s = {(lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = {lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2
      , (lut_in_data_sva_154[118:96])};
  wire[7:0] lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire[8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s = {(lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm[0]))};
  wire [48:0] nl_lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  wire [158:0] nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_else_else_le_index_u_1_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg_a;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0];
  wire [158:0] nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_1_lo_index_u_1_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  wire [158:0] nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_else_else_le_index_u_2_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg_a;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0];
  wire [158:0] nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_1_lo_index_u_2_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  wire [158:0] nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_else_else_le_index_u_3_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg_a;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0];
  wire [158:0] nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_1_lo_index_u_3_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  wire [158:0] nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_else_else_le_index_u_sva_3 , 127'b0};
  wire [48:0] nl_lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg_a;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0];
  wire [158:0] nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  assign nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a
      = {lut_lookup_else_1_lo_index_u_sva_3 , 127'b0};
  wire [323:0] nl_NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst_chn_lut_out_rsci_d;
  assign nl_NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst_chn_lut_out_rsci_d
      = {chn_lut_out_rsci_d_323 , chn_lut_out_rsci_d_322 , chn_lut_out_rsci_d_321
      , chn_lut_out_rsci_d_320 , chn_lut_out_rsci_d_319 , chn_lut_out_rsci_d_318
      , chn_lut_out_rsci_d_317 , chn_lut_out_rsci_d_316 , chn_lut_out_rsci_d_315
      , chn_lut_out_rsci_d_314 , chn_lut_out_rsci_d_313 , chn_lut_out_rsci_d_312_307
      , chn_lut_out_rsci_d_306 , chn_lut_out_rsci_d_305 , chn_lut_out_rsci_d_304
      , chn_lut_out_rsci_d_303_298 , chn_lut_out_rsci_d_297 , chn_lut_out_rsci_d_296
      , chn_lut_out_rsci_d_295 , chn_lut_out_rsci_d_294_289 , chn_lut_out_rsci_d_288
      , chn_lut_out_rsci_d_287 , chn_lut_out_rsci_d_286 , chn_lut_out_rsci_d_285_280
      , chn_lut_out_rsci_d_279 , chn_lut_out_rsci_d_278 , chn_lut_out_rsci_d_277
      , chn_lut_out_rsci_d_276 , chn_lut_out_rsci_d_275 , chn_lut_out_rsci_d_274
      , chn_lut_out_rsci_d_273 , chn_lut_out_rsci_d_272 , chn_lut_out_rsci_d_271
      , chn_lut_out_rsci_d_270 , chn_lut_out_rsci_d_269 , chn_lut_out_rsci_d_268
      , chn_lut_out_rsci_d_267_140 , chn_lut_out_rsci_d_139_117 , chn_lut_out_rsci_d_116_105
      , chn_lut_out_rsci_d_104_82 , chn_lut_out_rsci_d_81_70 , chn_lut_out_rsci_d_69_47
      , chn_lut_out_rsci_d_46_35 , chn_lut_out_rsci_d_34_12 , chn_lut_out_rsci_d_11_0};
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd32)) cfg_lut_le_start_rsci (
      .d(cfg_lut_le_start_rsci_d),
      .z(cfg_lut_le_start_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd32)) cfg_lut_lo_start_rsci (
      .d(cfg_lut_lo_start_rsci_d),
      .z(cfg_lut_lo_start_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd4),
  .width(32'sd8)) cfg_lut_le_index_offset_rsci (
      .d(cfg_lut_le_index_offset_rsci_d),
      .z(cfg_lut_le_index_offset_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd5),
  .width(32'sd8)) cfg_lut_le_index_select_rsci (
      .d(cfg_lut_le_index_select_rsci_d),
      .z(cfg_lut_le_index_select_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd6),
  .width(32'sd8)) cfg_lut_lo_index_select_rsci (
      .d(cfg_lut_lo_index_select_rsci_d),
      .z(cfg_lut_lo_index_select_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd7),
  .width(32'sd1)) cfg_lut_le_function_rsci (
      .d(cfg_lut_le_function_rsci_d),
      .z(cfg_lut_le_function_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd8),
  .width(32'sd1)) cfg_lut_uflow_priority_rsci (
      .d(cfg_lut_uflow_priority_rsci_d),
      .z(cfg_lut_uflow_priority_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd9),
  .width(32'sd1)) cfg_lut_oflow_priority_rsci (
      .d(cfg_lut_oflow_priority_rsci_d),
      .z(cfg_lut_oflow_priority_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd10),
  .width(32'sd1)) cfg_lut_hybrid_priority_rsci (
      .d(cfg_lut_hybrid_priority_rsci_d),
      .z(cfg_lut_hybrid_priority_rsc_z)
    );
  SDP_Y_IDX_mgc_in_wire_v1 #(.rscid(32'sd11),
  .width(32'sd2)) cfg_precision_rsci (
      .d(cfg_precision_rsci_d),
      .z(cfg_precision_rsc_z)
    );
  SDP_Y_IDX_leading_sign_32_0  lut_lookup_1_leading_sign_32_0_rg (
      .mantissa(lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0),
      .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_4)
    );
  SDP_Y_IDX_leading_sign_32_0  lut_lookup_2_leading_sign_32_0_rg (
      .mantissa(lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0),
      .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_5)
    );
  SDP_Y_IDX_leading_sign_32_0  lut_lookup_3_leading_sign_32_0_rg (
      .mantissa(lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0),
      .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_6)
    );
  SDP_Y_IDX_leading_sign_32_0  lut_lookup_4_leading_sign_32_0_rg (
      .mantissa(lut_lookup_if_else_else_le_data_sub_sva_mx0w0),
      .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_7)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg
      (
      .a(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
      .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg
      (
      .a(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
      .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg
      (
      .a(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s[8:0]),
      .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg
      (
      .a(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
      .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg
      (
      .a(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
      .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg
      (
      .a(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
      .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg
      (
      .a(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s[8:0]),
      .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg
      (
      .a(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
      .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg
      (
      .a(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
      .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg
      (
      .a(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
      .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg
      (
      .a(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s[8:0]),
      .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg
      (
      .a(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
      .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg
      (
      .a(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
      .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg
      (
      .a(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
      .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg
      (
      .a(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s[8:0]),
      .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd10),
  .width_z(32'sd256)) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg
      (
      .a(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a[23:0]),
      .s(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
      .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd35)) lut_lookup_1_if_else_else_else_else_if_lshift_rg (
      .a(nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_a[30:0]),
      .s(nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_s[5:0]),
      .z(lut_lookup_1_if_else_else_else_else_if_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd35)) lut_lookup_1_if_else_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_a[30:0]),
      .s(nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_s[7:0]),
      .z(lut_lookup_1_if_else_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_1_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_1_else_else_else_else_rshift_rg_a[34:0]),
      .s(nl_lut_lookup_1_else_else_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_1_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_1_else_1_else_else_rshift_rg (
      .a(lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2),
      .s(nl_lut_lookup_1_else_1_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_1_else_1_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd35)) lut_lookup_2_if_else_else_else_else_if_lshift_rg (
      .a(nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_a[30:0]),
      .s(nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_s[5:0]),
      .z(lut_lookup_2_if_else_else_else_else_if_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd35)) lut_lookup_2_if_else_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_a[30:0]),
      .s(nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_s[7:0]),
      .z(lut_lookup_2_if_else_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_2_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_2_else_else_else_else_rshift_rg_a[34:0]),
      .s(nl_lut_lookup_2_else_else_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_2_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_2_else_1_else_else_rshift_rg (
      .a(lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2),
      .s(nl_lut_lookup_2_else_1_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_2_else_1_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd35)) lut_lookup_3_if_else_else_else_else_if_lshift_rg (
      .a(nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_a[30:0]),
      .s(nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_s[5:0]),
      .z(lut_lookup_3_if_else_else_else_else_if_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd35)) lut_lookup_3_if_else_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_a[30:0]),
      .s(nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_s[7:0]),
      .z(lut_lookup_3_if_else_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_3_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_3_else_else_else_else_rshift_rg_a[34:0]),
      .s(nl_lut_lookup_3_else_else_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_3_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_3_else_1_else_else_rshift_rg (
      .a(lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2),
      .s(nl_lut_lookup_3_else_1_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_3_else_1_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd35)) lut_lookup_4_if_else_else_else_else_if_lshift_rg (
      .a(nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_a[30:0]),
      .s(nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_s[5:0]),
      .z(lut_lookup_4_if_else_else_else_else_if_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd31),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd35)) lut_lookup_4_if_else_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_a[30:0]),
      .s(nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_s[7:0]),
      .z(lut_lookup_4_if_else_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_4_else_else_else_else_rshift_rg (
      .a(nl_lut_lookup_4_else_else_else_else_rshift_rg_a[34:0]),
      .s(nl_lut_lookup_4_else_else_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_4_else_else_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd35)) lut_lookup_4_else_1_else_else_rshift_rg (
      .a(lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2),
      .s(nl_lut_lookup_4_else_1_else_else_rshift_rg_s[8:0]),
      .z(lut_lookup_4_else_1_else_else_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd32),
  .width_z(32'sd31)) lut_lookup_1_IntLog2_32U_lshift_rg (
      .a(1'b1),
      .s(nl_lut_lookup_1_IntLog2_32U_lshift_rg_s[31:0]),
      .z(lut_lookup_1_IntLog2_32U_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd32),
  .width_z(32'sd31)) lut_lookup_2_IntLog2_32U_lshift_rg (
      .a(1'b1),
      .s(nl_lut_lookup_2_IntLog2_32U_lshift_rg_s[31:0]),
      .z(lut_lookup_2_IntLog2_32U_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd32),
  .width_z(32'sd31)) lut_lookup_3_IntLog2_32U_lshift_rg (
      .a(1'b1),
      .s(nl_lut_lookup_3_IntLog2_32U_lshift_rg_s[31:0]),
      .z(lut_lookup_3_IntLog2_32U_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd32),
  .width_z(32'sd31)) lut_lookup_4_IntLog2_32U_lshift_rg (
      .a(1'b1),
      .s(nl_lut_lookup_4_IntLog2_32U_lshift_rg_s[31:0]),
      .z(lut_lookup_4_IntLog2_32U_lshift_itm)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_1_leading_sign_49_0_rg (
      .mantissa(nl_lut_lookup_1_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_1_leading_sign_49_0_2_rg (
      .mantissa(nl_lut_lookup_1_leading_sign_49_0_2_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_2_leading_sign_49_0_rg (
      .mantissa(nl_lut_lookup_2_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_2_leading_sign_49_0_2_rg (
      .mantissa(nl_lut_lookup_2_leading_sign_49_0_2_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_3_leading_sign_49_0_rg (
      .mantissa(nl_lut_lookup_3_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_3_leading_sign_49_0_2_rg (
      .mantissa(nl_lut_lookup_3_leading_sign_49_0_2_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_4_leading_sign_49_0_rg (
      .mantissa(nl_lut_lookup_4_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18)
    );
  SDP_Y_IDX_leading_sign_49_0  lut_lookup_4_leading_sign_49_0_2_rg (
      .mantissa(nl_lut_lookup_4_leading_sign_49_0_2_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_19_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_1_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_1_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_a_int_mant_p1_1_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_13_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_2_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_2_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_a_int_mant_p1_2_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_7_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_3_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_3_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_a_int_mant_p1_3_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_1_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_sva)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
      .a(nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_2_a_int_mant_p1_sva)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12),
      .z(lut_lookup_1_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_le_index_select_1_sva_5),
      .z(lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg (
      .a(nl_lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13),
      .z(lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_lo_index_select_1_sva_5),
      .z(lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14),
      .z(lut_lookup_2_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_le_index_select_1_sva_5),
      .z(lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg (
      .a(nl_lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15),
      .z(lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_lo_index_select_1_sva_5),
      .z(lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16),
      .z(lut_lookup_3_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_le_index_select_1_sva_5),
      .z(lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg (
      .a(nl_lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17),
      .z(lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_lo_index_select_1_sva_5),
      .z(lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18),
      .z(lut_lookup_4_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_le_index_select_1_sva_5),
      .z(lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg (
      .a(nl_lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19),
      .z(lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_itm)
    );
  SDP_Y_IDX_mgc_shift_br_v4 #(.width_a(32'sd159),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd287)) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg
      (
      .a(nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a[158:0]),
      .s(cfg_lut_lo_index_select_1_sva_5),
      .z(lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd32)) lut_lookup_1_else_else_else_else_le_data_f_lshift_1_rg (
      .a(1'b1),
      .s(cfg_lut_le_index_select_1_sva_6),
      .z(lut_lookup_1_else_else_else_else_le_data_f_lshift_1_itm)
    );
  SDP_Y_IDX_mgc_shift_bl_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd32)) lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_rg (
      .a(1'b1),
      .s(cfg_lut_lo_index_select_1_sva_6),
      .z(lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_itm)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_in_rsc_z(chn_lut_in_rsc_z),
      .chn_lut_in_rsc_vz(chn_lut_in_rsc_vz),
      .chn_lut_in_rsc_lz(chn_lut_in_rsc_lz),
      .chn_lut_in_rsci_oswt(chn_lut_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_lut_in_rsci_iswt0(chn_lut_in_rsci_iswt0),
      .chn_lut_in_rsci_bawt(chn_lut_in_rsci_bawt),
      .chn_lut_in_rsci_wen_comp(chn_lut_in_rsci_wen_comp),
      .chn_lut_in_rsci_ld_core_psct(chn_lut_in_rsci_ld_core_psct),
      .chn_lut_in_rsci_d_mxwt(chn_lut_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_out_rsc_z(chn_lut_out_rsc_z),
      .chn_lut_out_rsc_vz(chn_lut_out_rsc_vz),
      .chn_lut_out_rsc_lz(chn_lut_out_rsc_lz),
      .chn_lut_out_rsci_oswt(chn_lut_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_lut_out_rsci_iswt0(chn_lut_out_rsci_iswt0),
      .chn_lut_out_rsci_bawt(chn_lut_out_rsci_bawt),
      .chn_lut_out_rsci_wen_comp(chn_lut_out_rsci_wen_comp),
      .chn_lut_out_rsci_ld_core_psct(reg_chn_lut_out_rsci_ld_core_psct_cse),
      .chn_lut_out_rsci_d(nl_NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst_chn_lut_out_rsci_d[323:0])
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_staller NV_NVDLA_SDP_CORE_Y_idx_core_staller_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_lut_in_rsci_wen_comp(chn_lut_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_lut_out_rsci_wen_comp(chn_lut_out_rsci_wen_comp)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign chn_lut_out_and_cse = core_wen & (~(and_dcpl_54 | (~ main_stage_v_5)));
  assign chn_lut_out_and_13_cse = core_wen & ((or_cse & main_stage_v_5 & lut_lookup_1_and_svs_2)
      | and_dcpl_59);
  assign chn_lut_out_and_14_cse = core_wen & ((or_cse & main_stage_v_5 & lut_lookup_2_and_svs_2)
      | and_dcpl_63);
  assign chn_lut_out_and_15_cse = core_wen & ((or_cse & main_stage_v_5 & lut_lookup_3_and_svs_2)
      | and_dcpl_67);
  assign chn_lut_out_and_16_cse = core_wen & ((or_cse & main_stage_v_5 & lut_lookup_4_and_svs_2)
      | and_dcpl_71);
  assign lut_lookup_and_138_cse = (~ lut_lookup_unequal_tmp_13) & lut_lookup_or_3_tmp;
  assign lut_lookup_and_139_cse = lut_lookup_unequal_tmp_13 & lut_lookup_or_3_tmp;
  assign lut_lookup_and_136_cse = (~ lut_lookup_unequal_tmp_13) & lut_lookup_or_7_tmp;
  assign lut_lookup_and_137_cse = lut_lookup_unequal_tmp_13 & lut_lookup_or_7_tmp;
  assign lut_lookup_and_134_cse = (~ lut_lookup_unequal_tmp_13) & lut_lookup_or_11_tmp;
  assign lut_lookup_and_135_cse = lut_lookup_unequal_tmp_13 & lut_lookup_or_11_tmp;
  assign lut_lookup_and_132_cse = (~ lut_lookup_unequal_tmp_13) & lut_lookup_or_15_tmp;
  assign lut_lookup_and_133_cse = lut_lookup_unequal_tmp_13 & lut_lookup_or_15_tmp;
  assign cfg_precision_and_cse = core_wen & (~ and_dcpl_54) & mux_580_cse;
  assign mux_4_nl = MUX_s_1_2_2(or_tmp_8, or_tmp_6, or_cse);
  assign FpAdd_8U_23U_2_is_addition_and_cse = core_wen & (~ and_dcpl_54) & (~ (mux_4_nl));
  assign FpAdd_8U_23U_1_is_addition_and_1_cse = core_wen & (~ and_dcpl_54) & (~ mux_tmp_4);
  assign cfg_lut_le_index_offset_and_1_cse = core_wen & (~ and_dcpl_54) & mux_tmp_10;
  assign or_26_cse = (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10);
  assign nor_783_nl = ~(or_cse | (~ or_66_cse));
  assign mux_1120_nl = MUX_s_1_2_2(or_tmp_1490, (nor_783_nl), reg_cfg_precision_1_sva_st_12_cse_1[1]);
  assign mux_1121_nl = MUX_s_1_2_2((mux_1120_nl), or_tmp_1490, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign FpAdd_8U_23U_1_mux1h_1_itm = MUX_v_8_2_2(FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5,
      ({2'b0 , libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_4}),
      mux_1121_nl);
  assign or_cse = chn_lut_out_rsci_bawt | (~ reg_chn_lut_out_rsci_ld_core_psct_cse);
  assign and_956_cse = (reg_cfg_precision_1_sva_st_12_cse_1==2'b10);
  assign and_284_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & (~ reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse);
  assign and_286_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_288_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse) & (~
      reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse);
  assign and_290_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse) & reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_2_and_35_cse = core_wen & (~ and_dcpl_54) & (~ mux_20_itm);
  assign and_292_rgt = or_cse & reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign mux_1122_cse = MUX_s_1_2_2(or_66_cse, or_26_cse, or_cse);
  assign FpAdd_8U_23U_1_mux1h_3_itm = MUX_v_8_2_2(FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5,
      ({2'b0 , libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_5}),
      mux_1122_cse);
  assign nor_874_cse = ~(chn_lut_out_rsci_bawt | (~ reg_chn_lut_out_rsci_ld_core_psct_cse));
  assign and_961_cse = and_dcpl_540 & (reg_cfg_precision_1_sva_st_12_cse_1[1]) &
      (~(nor_874_cse | (reg_cfg_precision_1_sva_st_12_cse_1[0])));
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse = (or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse)
      | and_524_rgt;
  assign IsNaN_8U_23U_3_aelse_and_3_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse
      & (~ mux_25_itm);
  assign and_300_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & (~ reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse);
  assign and_302_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_304_rgt = or_cse & (~(reg_cfg_lut_le_function_1_sva_st_19_cse | reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse));
  assign and_306_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse) & reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_2_and_36_cse = core_wen & (~ and_dcpl_54) & (~ mux_26_itm);
  assign and_308_rgt = or_cse & reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_1_mux1h_5_itm = MUX_v_8_2_2(FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5,
      ({2'b0 , libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_6}),
      mux_1122_cse);
  assign and_316_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & (~ reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse);
  assign and_318_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_320_rgt = or_cse & (~(reg_cfg_lut_le_function_1_sva_st_19_cse | reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse));
  assign and_322_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse) & reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_2_and_37_cse = core_wen & (~ and_dcpl_54) & (~ mux_25_itm);
  assign and_324_rgt = or_cse & reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_1_mux1h_7_itm = MUX_v_8_2_2(FpAdd_8U_23U_1_qr_lpi_1_dfm_5,
      ({2'b0 , libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_7}),
      mux_1122_cse);
  assign and_330_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & (~ reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse);
  assign and_332_rgt = or_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_334_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse) & (~
      reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse);
  assign and_336_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse) & reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_338_rgt = or_cse & reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign cfg_lut_le_start_and_cse = core_wen & (~ and_dcpl_54) & mux_tmp_35;
  assign and_344_rgt = (~ or_66_cse) & (~ reg_cfg_lut_le_function_1_sva_st_20_cse)
      & or_cse;
  assign and_347_rgt = or_66_cse & (~ reg_cfg_lut_le_function_1_sva_st_20_cse) &
      or_cse;
  assign or_66_cse = (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10);
  assign nor_792_cse = ~((cfg_precision_1_sva_st_70!=2'b10));
  assign nor_775_nl = ~(nor_5_cse_1 | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 | IsNaN_8U_23U_4_land_1_lpi_1_dfm_4
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10));
  assign nor_776_nl = ~(IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 |
      (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign mux_42_nl = MUX_s_1_2_2((nor_776_nl), (nor_775_nl), or_cse);
  assign FpMantRNE_49U_24U_1_else_o_mant_and_cse = core_wen & (~ and_dcpl_54) & (mux_42_nl);
  assign and_355_m1c = or_dcpl_51 & or_cse;
  assign nor_5_cse_1 = ~(lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 | (~ (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49])));
  assign nl_lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm}) + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)})
      + 8'b1;
  assign lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt = nl_lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt[7:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm}) + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt = nl_lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt[7:0];
  assign FpAdd_8U_23U_o_expo_and_3_ssc = (~ (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]))
      & and_355_m1c;
  assign FpAdd_8U_23U_and_51_ssc = (~ lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7)
      & (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]) & and_355_m1c;
  assign FpAdd_8U_23U_and_43_ssc = lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7
      & (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]) & and_355_m1c;
  assign mux_1220_nl = MUX_s_1_2_2(IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5, IsNaN_8U_23U_4_land_1_lpi_1_dfm_4,
      reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign or_1936_cse = (~((mux_1220_nl) | nor_5_cse_1 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_7))
      | lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
  assign nor_865_cse = ~(nor_874_cse | (reg_cfg_precision_1_sva_st_13_cse_1[0]));
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse = ((~ or_66_cse) & or_cse) | and_dcpl_161;
  assign IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse = and_dcpl_148 | and_dcpl_162;
  assign IsNaN_8U_23U_3_aelse_and_6_cse = core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse
      & (~ mux_83_cse);
  assign FpMantRNE_49U_24U_1_else_and_cse = core_wen & (~ and_dcpl_54) & (~ mux_83_cse);
  assign nor_13_cse = ~(lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49])));
  assign FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse =
      and_401_cse | and_dcpl_161;
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt = ~((FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49])
      | and_dcpl_54);
  assign FpAdd_8U_23U_2_and_4_rgt = (~ lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49]) & (~ and_dcpl_54);
  assign FpAdd_8U_23U_2_and_5_rgt = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49]) & (~ and_dcpl_54);
  assign mux_83_cse = MUX_s_1_2_2(or_tmp_63, or_1689_cse, or_cse);
  assign FpAdd_8U_23U_2_is_inf_and_cse = core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
      & mux_tmp_35;
  assign and_364_rgt = and_dcpl_98 & (~ reg_cfg_lut_le_function_1_sva_st_20_cse)
      & or_cse;
  assign IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse = and_364_rgt | and_dcpl_148
      | and_347_rgt;
  assign nor_764_nl = ~(nor_27_cse_1 | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10)
      | IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_4_land_2_lpi_1_dfm_5);
  assign nor_765_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10) |
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6
      | FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6);
  assign mux_92_nl = MUX_s_1_2_2((nor_765_nl), (nor_764_nl), or_cse);
  assign FpMantRNE_49U_24U_1_else_o_mant_and_1_cse = core_wen & (~ and_dcpl_54) &
      (mux_92_nl);
  assign and_375_m1c = or_dcpl_57 & or_cse;
  assign nor_27_cse_1 = ~(lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 | (~ (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49])));
  assign nl_lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm}) + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)})
      + 8'b1;
  assign lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt = nl_lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt[7:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm}) + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt = nl_lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt[7:0];
  assign FpAdd_8U_23U_o_expo_and_2_ssc = (~ (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]))
      & and_375_m1c;
  assign FpAdd_8U_23U_and_53_ssc = (~ lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7)
      & (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]) & and_375_m1c;
  assign FpAdd_8U_23U_and_45_ssc = lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7
      & (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]) & and_375_m1c;
  assign mux_1227_nl = MUX_s_1_2_2(IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5, IsNaN_8U_23U_4_land_2_lpi_1_dfm_5,
      reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign nor_855_cse = ~((mux_1227_nl) | nor_27_cse_1 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_7);
  assign mux_1126_cse = MUX_s_1_2_2(and_896_cse, or_dcpl_57, or_cse);
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse = (and_dcpl_98 & or_cse) | and_dcpl_161;
  assign FpAdd_8U_23U_1_is_inf_and_1_cse = core_wen & FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse
      & mux_tmp_35;
  assign nor_31_cse = ~(lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49])));
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt = ~((FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49])
      | and_dcpl_54);
  assign FpAdd_8U_23U_2_and_10_rgt = (~ lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49]) & (~ and_dcpl_54);
  assign FpAdd_8U_23U_2_and_11_rgt = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49]) & (~ and_dcpl_54);
  assign mux_132_nl = MUX_s_1_2_2(or_tmp_63, or_tmp_44, or_cse);
  assign IsNaN_8U_23U_8_aelse_and_1_cse = core_wen & (~ and_dcpl_54) & (~ (mux_132_nl));
  assign or_48_cse = (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7) | reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign nor_749_nl = ~(nor_38_cse_1 | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10)
      | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      | IsNaN_8U_23U_4_land_3_lpi_1_dfm_5);
  assign nor_750_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10) |
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6
      | FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6);
  assign mux_141_nl = MUX_s_1_2_2((nor_750_nl), (nor_749_nl), or_cse);
  assign FpMantRNE_49U_24U_1_else_o_mant_and_2_cse = core_wen & (~ and_dcpl_54) &
      (mux_141_nl);
  assign nor_38_cse_1 = ~(lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 | (~ (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49])));
  assign nl_lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm}) + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16)})
      + 8'b1;
  assign lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt = nl_lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt[7:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm}) + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt = nl_lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt[7:0];
  assign FpAdd_8U_23U_o_expo_and_1_ssc = (~ (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]))
      & and_375_m1c;
  assign FpAdd_8U_23U_and_55_ssc = (~ lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7)
      & (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]) & and_375_m1c;
  assign FpAdd_8U_23U_and_47_ssc = lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7
      & (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]) & and_375_m1c;
  assign nor_42_cse = ~(lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49])));
  assign and_401_cse = (reg_cfg_precision_1_sva_st_13_cse_1==2'b10) & or_cse;
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt = ~((FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49])
      | and_dcpl_54);
  assign FpAdd_8U_23U_2_and_16_rgt = (~ lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49]) & (~ and_dcpl_54);
  assign FpAdd_8U_23U_2_and_17_rgt = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49]) & (~ and_dcpl_54);
  assign nor_737_nl = ~(nor_50_cse_1 | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10)
      | reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse | IsNaN_8U_23U_1_land_lpi_1_dfm_7
      | IsNaN_8U_23U_4_land_lpi_1_dfm_4);
  assign nor_738_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10) |
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 | IsNaN_8U_23U_3_land_lpi_1_dfm_6 | IsNaN_8U_23U_3_land_lpi_1_dfm_st_6
      | FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6);
  assign mux_177_nl = MUX_s_1_2_2((nor_738_nl), (nor_737_nl), or_cse);
  assign FpMantRNE_49U_24U_1_else_o_mant_and_3_cse = core_wen & (~ and_dcpl_54) &
      (mux_177_nl);
  assign nor_50_cse_1 = ~(lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 | (~ (FpAdd_8U_23U_1_int_mant_p1_sva_3[49])));
  assign nl_lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm}) + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18)})
      + 8'b1;
  assign lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt = nl_lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt[7:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt = ({reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm
      , reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm}) + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt = nl_lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt[7:0];
  assign FpAdd_8U_23U_o_expo_and_ssc = (~ (FpAdd_8U_23U_1_int_mant_p1_sva_3[49]))
      & and_375_m1c;
  assign FpAdd_8U_23U_and_57_ssc = (~ lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7)
      & (FpAdd_8U_23U_1_int_mant_p1_sva_3[49]) & and_375_m1c;
  assign FpAdd_8U_23U_and_49_ssc = lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7
      & (FpAdd_8U_23U_1_int_mant_p1_sva_3[49]) & and_375_m1c;
  assign nor_54_cse = ~(lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_2_int_mant_p1_sva_3[49])));
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt = ~((FpAdd_8U_23U_2_int_mant_p1_sva_3[49])
      | and_dcpl_54);
  assign FpAdd_8U_23U_2_and_22_rgt = (~ lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_2_int_mant_p1_sva_3[49]) & (~ and_dcpl_54);
  assign FpAdd_8U_23U_2_and_23_rgt = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_2_int_mant_p1_sva_3[49]) & (~ and_dcpl_54);
  assign and_428_rgt = and_896_cse & or_cse;
  assign and_427_cse = or_1857_cse & or_cse;
  assign or_312_cse = (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse
      = and_427_cse | and_428_rgt;
  assign nor_724_nl = ~(cfg_lut_le_function_1_sva_st_41 | (~ and_tmp_6));
  assign nor_725_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~(main_stage_v_4 & or_tmp_314)));
  assign mux_220_nl = MUX_s_1_2_2((nor_725_nl), (nor_724_nl), or_cse);
  assign lut_lookup_if_else_if_and_cse = core_wen & (~ and_dcpl_54) & (mux_220_nl);
  assign cfg_precision_and_24_cse = core_wen & (~ and_dcpl_54) & mux_tmp_220;
  assign nor_722_nl = ~((~ cfg_lut_le_function_1_sva_st_41) | and_1142_cse | FpAdd_8U_23U_1_mux_13_itm_4
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp | (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign nor_723_nl = ~((~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign mux_222_nl = MUX_s_1_2_2((nor_723_nl), (nor_722_nl), or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse = core_wen & (~ and_dcpl_54)
      & (mux_222_nl);
  assign and_430_rgt = or_cse & (~ cfg_lut_le_function_1_sva_st_41);
  assign FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse = (or_cse & cfg_lut_le_function_1_sva_st_41)
      | and_430_rgt;
  assign or_332_nl = lut_lookup_if_1_lor_5_lpi_1_dfm_4 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_226_nl = MUX_s_1_2_2((or_332_nl), or_tmp_331, or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse = core_wen & (~ and_dcpl_54)
      & (~ (mux_226_nl));
  assign nor_715_nl = ~((~ cfg_lut_le_function_1_sva_st_41) | IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp | FpAdd_8U_23U_1_mux_29_itm_4 |
      (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign nor_716_nl = ~((~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign mux_234_nl = MUX_s_1_2_2((nor_716_nl), (nor_715_nl), or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse = core_wen & (~ and_dcpl_54)
      & (mux_234_nl);
  assign or_365_cse = lut_lookup_if_1_lor_6_lpi_1_dfm_4 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_238_nl = MUX_s_1_2_2(or_365_cse, or_tmp_363, or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse = core_wen & (~ and_dcpl_54)
      & (~ (mux_238_nl));
  assign or_1857_cse = (cfg_precision_1_sva_st_70!=2'b10);
  assign nor_707_nl = ~((~ cfg_lut_le_function_1_sva_st_41) | IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp | FpAdd_8U_23U_1_mux_45_itm_4 |
      (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign nor_708_nl = ~((~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign mux_247_nl = MUX_s_1_2_2((nor_708_nl), (nor_707_nl), or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse = core_wen & (~ and_dcpl_54)
      & (mux_247_nl);
  assign mux_251_nl = MUX_s_1_2_2(or_tmp_397, or_tmp_395, or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse = core_wen & (~ and_dcpl_54)
      & (~ (mux_251_nl));
  assign nor_701_nl = ~((~ cfg_lut_le_function_1_sva_st_41) | IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp | FpAdd_8U_23U_1_mux_61_itm_4
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign nor_702_nl = ~((~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign mux_259_nl = MUX_s_1_2_2((nor_702_nl), (nor_701_nl), or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse = core_wen & (~ and_dcpl_54)
      & (mux_259_nl);
  assign mux_263_nl = MUX_s_1_2_2(or_tmp_428, or_tmp_427, or_cse);
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse = core_wen & (~ and_dcpl_54)
      & (~ (mux_263_nl));
  assign cfg_lut_hybrid_priority_and_cse = core_wen & (~ and_dcpl_54) & mux_tmp_265;
  assign lut_lookup_else_mux_180_cse = MUX_s_1_2_2(lut_lookup_if_mux_mx0w1, lut_lookup_else_mux_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign or_1853_cse = (~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_else_unequal_tmp_18;
  assign and_854_cse = or_1853_cse & lut_lookup_else_if_lor_5_lpi_1_dfm_5;
  assign mux_275_nl = MUX_s_1_2_2(or_tmp_456, or_tmp_380, or_cse);
  assign lut_lookup_else_if_oelse_1_and_1_cse = core_wen & (~ and_dcpl_54) & (~ (mux_275_nl));
  assign and_852_cse = cfg_lut_le_function_1_sva_st_42 & main_stage_v_4;
  assign nor_690_cse = ~(lut_lookup_if_1_lor_5_lpi_1_dfm_4 | (~ main_stage_v_4) |
      (cfg_precision_1_sva_st_71!=2'b10));
  assign and_846_cse = lut_lookup_unequal_tmp_13 & lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  assign mux_283_cse = MUX_s_1_2_2((~ main_stage_v_5), or_tmp_478, lut_lookup_unequal_tmp_13);
  assign mux_284_nl = MUX_s_1_2_2(mux_283_cse, mux_tmp_281, or_cse);
  assign lut_lookup_if_1_oelse_1_and_4_cse = core_wen & (~ and_dcpl_54) & (~ (mux_284_nl));
  assign mux_285_nl = MUX_s_1_2_2(or_tmp_478, or_312_cse, or_cse);
  assign lut_lookup_if_1_oelse_1_and_5_cse = core_wen & (~ and_dcpl_54) & (~ (mux_285_nl));
  assign lut_lookup_else_mux_182_cse = MUX_s_1_2_2(lut_lookup_if_mux_41_mx0w1, lut_lookup_else_mux_43_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign or_492_cse = (~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_else_unequal_tmp_12;
  assign and_82_cse = lut_lookup_else_if_lor_6_lpi_1_dfm_5 & or_492_cse;
  assign and_843_cse = cfg_lut_le_function_1_sva_10 & main_stage_v_5;
  assign lut_lookup_else_mux_184_cse = MUX_s_1_2_2(lut_lookup_if_mux_82_mx0w1, lut_lookup_else_mux_86_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign and_839_cse = or_492_cse & lut_lookup_else_if_lor_7_lpi_1_dfm_5;
  assign mux_314_nl = MUX_s_1_2_2(or_tmp_456, (~ main_stage_v_5), cfg_lut_le_function_1_sva_10);
  assign mux_315_nl = MUX_s_1_2_2((mux_314_nl), or_tmp_456, lut_lookup_else_unequal_tmp_13);
  assign mux_316_nl = MUX_s_1_2_2((mux_315_nl), mux_tmp_292, or_cse);
  assign lut_lookup_else_if_oelse_1_and_4_cse = core_wen & (~ and_dcpl_54) & (~ (mux_316_nl));
  assign mux_328_nl = MUX_s_1_2_2(mux_283_cse, or_312_cse, or_cse);
  assign mux_329_nl = MUX_s_1_2_2(mux_283_cse, (~ main_stage_v_4), or_cse);
  assign mux_330_nl = MUX_s_1_2_2((mux_329_nl), (mux_328_nl), lut_lookup_else_unequal_tmp_18);
  assign lut_lookup_if_1_oelse_1_and_8_cse = core_wen & (~ and_dcpl_54) & (~ (mux_330_nl));
  assign lut_lookup_else_mux_186_cse = MUX_s_1_2_2(lut_lookup_if_mux_123_mx0w1, lut_lookup_else_mux_129_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign and_835_cse = or_492_cse & lut_lookup_else_if_lor_1_lpi_1_dfm_5;
  assign lut_lookup_le_uflow_and_cse = core_wen & (and_dcpl_258 | and_dcpl_259) &
      mux_tmp_265;
  assign mux_356_nl = MUX_s_1_2_2(and_832_cse, main_stage_v_4, or_cse);
  assign nor_657_nl = ~((~ reg_chn_lut_out_rsci_ld_core_psct_cse) | chn_lut_out_rsci_bawt
      | (~ and_832_cse));
  assign mux_357_nl = MUX_s_1_2_2((nor_657_nl), (mux_356_nl), lut_lookup_else_unequal_tmp_18);
  assign lut_lookup_lo_index_0_and_cse = core_wen & (~ and_dcpl_54) & (mux_357_nl);
  assign and_465_cse = or_1202_cse & and_dcpl_259;
  assign and_466_cse = (~ or_1202_cse) & and_dcpl_259;
  assign lut_lookup_else_else_lut_lookup_else_else_or_3_cse = and_dcpl_258 | and_465_cse
      | and_466_cse;
  assign mux_358_nl = MUX_s_1_2_2(nor_612_cse, main_stage_v_4, lut_lookup_else_unequal_tmp_12);
  assign mux_359_nl = MUX_s_1_2_2(not_tmp_334, main_stage_v_5, lut_lookup_else_unequal_tmp_13);
  assign mux_360_nl = MUX_s_1_2_2((mux_359_nl), (mux_358_nl), or_cse);
  assign lut_lookup_else_else_and_cse = core_wen & lut_lookup_else_else_lut_lookup_else_else_or_3_cse
      & (mux_360_nl);
  assign and_832_cse = lut_lookup_unequal_tmp_13 & main_stage_v_5;
  assign mux_366_nl = MUX_s_1_2_2(and_832_cse, nor_tmp_112, or_cse);
  assign lut_lookup_lo_index_0_and_2_cse = core_wen & (~ and_dcpl_54) & (mux_366_nl);
  assign lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse = and_427_cse | and_636_cse;
  assign lut_lookup_lo_uflow_and_4_cse = core_wen & lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse
      & mux_tmp_220;
  assign lut_lookup_FpAdd_8U_23U_1_or_11_cse = (FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse
      & or_cse) | and_dcpl_280;
  assign FpAdd_8U_23U_1_and_46_cse = core_wen & lut_lookup_FpAdd_8U_23U_1_or_11_cse
      & (~ mux_3_itm);
  assign lut_lookup_FpAdd_8U_23U_2_or_10_cse = (FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse
      & or_cse) | and_dcpl_292;
  assign FpAdd_8U_23U_2_and_44_cse = core_wen & lut_lookup_FpAdd_8U_23U_2_or_10_cse
      & (~ mux_tmp_4);
  assign lut_lookup_FpAdd_8U_23U_2_or_9_cse = (FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse
      & or_cse) | and_dcpl_300;
  assign lut_lookup_FpAdd_8U_23U_2_or_8_cse = (FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse
      & or_cse) | and_dcpl_308;
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1)
      & lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_4_itm_8_1;
  assign FpAdd_8U_23U_1_is_a_greater_oelse_and_cse = core_wen & ((and_dcpl_309 &
      cfg_lut_le_function_rsci_d & or_cse) | (and_dcpl_309 & (~ cfg_lut_le_function_rsci_d)
      & or_cse) | and_dcpl_314) & mux_580_cse;
  assign IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse = and_dcpl_315 | and_dcpl_316;
  assign IsZero_8U_23U_4_and_cse = core_wen & IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse
      & (~ mux_3_itm);
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse = ((~ FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_itm_23_1)
      & lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_2_is_a_greater_acc_itm_8_1;
  assign FpAdd_8U_23U_2_is_a_greater_oelse_and_cse = core_wen & ((and_dcpl_309 &
      or_cse) | and_dcpl_314) & mux_580_cse;
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1)
      & lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_6_itm_8_1;
  assign IsZero_8U_23U_4_and_1_cse = core_wen & IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse
      & (~ mux_tmp_4);
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse = ((~ FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_itm_23_1)
      & lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_2_is_a_greater_acc_1_itm_8_1;
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1)
      & lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_8_itm_8_1;
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse = ((~ FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_itm_23_1)
      & lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_2_is_a_greater_acc_2_itm_8_1;
  assign mux_580_cse = MUX_s_1_2_2(main_stage_v_1, chn_lut_in_rsci_bawt, or_cse);
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1)
      & lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_10_itm_8_1;
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse = ((~ FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_itm_23_1)
      & lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_2_is_a_greater_acc_3_itm_8_1;
  assign IsZero_8U_23U_7_and_3_cse = core_wen & (~ and_dcpl_54) & (~ mux_595_itm);
  assign and_524_rgt = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse);
  assign and_525_rgt = or_26_cse & or_cse;
  assign IsNaN_8U_23U_1_aelse_and_4_cse = core_wen & (((reg_cfg_precision_1_sva_st_12_cse_1==2'b10)
      & or_cse) | and_525_rgt) & mux_tmp_10;
  assign and_527_rgt = and_956_cse & (~ reg_cfg_lut_le_function_1_sva_st_19_cse)
      & or_cse;
  assign and_529_rgt = and_956_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & or_cse;
  assign IsNaN_8U_23U_1_aelse_and_5_cse = core_wen & (and_527_rgt | and_529_rgt |
      and_525_rgt) & mux_tmp_10;
  assign IsNaN_8U_23U_7_aelse_and_17_cse = core_wen & ((and_956_cse & or_cse) | and_525_rgt)
      & mux_tmp_10;
  assign mux_1185_nl = MUX_s_1_2_2(IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4, IsNaN_8U_23U_1_land_1_lpi_1_dfm_6,
      reg_cfg_lut_le_function_1_sva_st_19_cse);
  assign and_551_rgt = (mux_1185_nl) & or_cse;
  assign lut_lookup_or_17_rgt = ((~ IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0) & and_553_m1c)
      | ((~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_6) & and_555_m1c);
  assign lut_lookup_or_18_rgt = (IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0 & and_553_m1c)
      | (IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 & and_555_m1c);
  assign and_562_m1c = main_stage_v_1 & (~ IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4)
      & (reg_cfg_precision_1_sva_st_12_cse_1[1]) & and_dcpl_351;
  assign nor_648_cse = ~((~ chn_lut_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10));
  assign or_1689_cse = (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10);
  assign and_559_rgt = main_stage_v_1 & IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 & (reg_cfg_precision_1_sva_st_12_cse_1[1])
      & and_dcpl_351;
  assign lut_lookup_and_126_rgt = (~ IsNaN_8U_23U_8_land_2_lpi_1_dfm_5) & and_562_m1c;
  assign lut_lookup_and_127_rgt = IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 & and_562_m1c;
  assign or_1688_cse = (~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10);
  assign and_564_rgt = or_1688_cse & main_stage_v_2 & and_401_cse;
  assign nor_190_cse = ~((reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign and_567_m1c = or_cse & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4);
  assign and_566_rgt = or_cse & IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign lut_lookup_and_124_rgt = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_6) & and_567_m1c;
  assign lut_lookup_and_125_rgt = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 & and_567_m1c;
  assign and_572_m1c = and_dcpl_364 & or_cse & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4);
  assign and_570_rgt = and_dcpl_364 & or_cse & IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign lut_lookup_and_122_rgt = (~ IsNaN_8U_23U_8_land_2_lpi_1_dfm_5) & and_572_m1c;
  assign lut_lookup_and_123_rgt = IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 & and_572_m1c;
  assign or_1691_cse = or_26_cse | (~ main_stage_v_1);
  assign and_574_rgt = or_1691_cse & main_stage_v_2 & and_401_cse;
  assign nor_193_cse = ~((reg_cfg_precision_1_sva_st_13_cse_1!=2'b10));
  assign and_577_m1c = or_cse & (~ IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4);
  assign and_576_rgt = or_cse & IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign lut_lookup_and_120_rgt = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_6) & and_577_m1c;
  assign lut_lookup_and_121_rgt = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 & and_577_m1c;
  assign and_582_m1c = and_dcpl_364 & or_cse & (~ IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4);
  assign and_580_rgt = and_dcpl_364 & or_cse & IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign lut_lookup_and_118_rgt = (~ nor_482_cse) & and_582_m1c;
  assign lut_lookup_and_119_rgt = nor_482_cse & and_582_m1c;
  assign and_586_rgt = or_1691_cse & (reg_cfg_precision_1_sva_st_13_cse_1==2'b10)
      & main_stage_v_2 & or_cse;
  assign or_849_cse = (~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign nor_196_cse = ~((~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign or_1696_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_6 | (~ reg_cfg_lut_le_function_1_sva_st_19_cse);
  assign and_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_6 & reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign mux_1186_nl = MUX_s_1_2_2((and_nl), (or_1696_nl), reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse);
  assign and_588_rgt = (mux_1186_nl) & or_cse;
  assign lut_lookup_or_rgt = ((~ IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0) & and_590_m1c)
      | ((~ IsNaN_8U_23U_1_land_lpi_1_dfm_6) & and_592_m1c);
  assign lut_lookup_or_16_rgt = (IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0 & and_590_m1c)
      | (IsNaN_8U_23U_1_land_lpi_1_dfm_6 & and_592_m1c);
  assign and_597_m1c = and_dcpl_364 & or_cse & (~ reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse);
  assign and_595_rgt = and_dcpl_364 & or_cse & reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign lut_lookup_and_112_rgt = (~ nor_469_cse) & and_597_m1c;
  assign lut_lookup_and_113_rgt = nor_469_cse & and_597_m1c;
  assign and_604_rgt = and_896_cse & cfg_lut_le_function_1_sva_st_41 & or_cse;
  assign and_606_rgt = or_1857_cse & (~ cfg_lut_le_function_1_sva_st_41) & or_cse;
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse = and_604_rgt | and_606_rgt
      | and_dcpl_403 | and_dcpl_405;
  assign mux_668_nl = MUX_s_1_2_2(or_tmp_63, (~ main_stage_v_3), cfg_precision_1_sva_st_70[1]);
  assign mux_1285_cse = MUX_s_1_2_2((mux_668_nl), or_tmp_63, cfg_precision_1_sva_st_70[0]);
  assign mux_670_cse = mux_1285_cse | (~ cfg_lut_le_function_1_sva_st_41);
  assign mux_671_nl = MUX_s_1_2_2(mux_tmp_292, mux_670_cse, or_cse);
  assign lut_lookup_else_if_oelse_1_and_8_cse = core_wen & (~ and_dcpl_54) & (~ (mux_671_nl));
  assign and_826_cse = cfg_lut_le_function_1_sva_st_41 & main_stage_v_3;
  assign nor_634_cse = ~((~ lut_lookup_else_unequal_tmp_12) | (cfg_precision_1_sva_st_71!=2'b10));
  assign mux_706_nl = MUX_s_1_2_2(main_stage_v_4, mux_tmp_704, or_cse);
  assign and_120_nl = or_cse & mux_tmp_704;
  assign mux_707_nl = MUX_s_1_2_2((and_120_nl), (mux_706_nl), lut_lookup_else_unequal_tmp_18);
  assign lut_lookup_lo_index_0_and_4_cse = core_wen & (~ and_dcpl_54) & (mux_707_nl);
  assign and_636_cse = (cfg_precision_1_sva_st_70==2'b10) & or_cse;
  assign mux_715_nl = MUX_s_1_2_2(or_312_cse, mux_1285_cse, or_cse);
  assign mux_716_nl = MUX_s_1_2_2((~ main_stage_v_4), mux_1285_cse, or_cse);
  assign mux_717_nl = MUX_s_1_2_2((mux_716_nl), (mux_715_nl), lut_lookup_else_unequal_tmp_18);
  assign lut_lookup_if_1_oelse_1_and_12_cse = core_wen & (~ and_dcpl_54) & (~ (mux_717_nl));
  assign mux_729_nl = MUX_s_1_2_2(nor_tmp_112, mux_tmp_704, or_cse);
  assign lut_lookup_lo_index_0_and_6_cse = core_wen & (~ and_dcpl_54) & (mux_729_nl);
  assign mux_735_nl = MUX_s_1_2_2(mux_tmp_281, mux_1285_cse, or_cse);
  assign lut_lookup_if_1_oelse_1_and_14_cse = core_wen & (~ and_dcpl_54) & (~ (mux_735_nl));
  assign or_969_cse = FpAdd_8U_23U_2_mux_13_itm_3 | and_1141_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp;
  assign or_978_cse = cfg_lut_le_function_1_sva_st_42 | (~ main_stage_v_4);
  assign mux_743_nl = MUX_s_1_2_2(or_tmp_976, (~ main_stage_v_3), cfg_precision_1_sva_st_70[1]);
  assign mux_1282_nl = MUX_s_1_2_2((mux_743_nl), or_tmp_976, cfg_precision_1_sva_st_70[0]);
  assign mux_745_cse = (mux_1282_nl) | cfg_lut_le_function_1_sva_st_41;
  assign mux_746_nl = MUX_s_1_2_2(or_tmp_980, (~ main_stage_v_4), cfg_precision_1_sva_st_71[1]);
  assign mux_747_nl = MUX_s_1_2_2((mux_746_nl), or_tmp_980, cfg_precision_1_sva_st_71[0]);
  assign mux_748_nl = MUX_s_1_2_2((mux_747_nl), or_978_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_749_nl = MUX_s_1_2_2((mux_748_nl), mux_745_cse, or_cse);
  assign lut_lookup_if_if_oelse_1_and_cse = core_wen & (~ and_dcpl_54) & (~ (mux_749_nl));
  assign mux_754_nl = MUX_s_1_2_2(main_stage_v_4, (~ or_tmp_993), cfg_precision_1_sva_st_71[1]);
  assign mux_755_cse = MUX_s_1_2_2((mux_754_nl), main_stage_v_4, cfg_precision_1_sva_st_71[0]);
  assign nor_612_cse = ~(cfg_lut_le_function_1_sva_st_42 | (~ main_stage_v_4));
  assign nor_610_cse = ~((cfg_precision_1_sva_8!=2'b10));
  assign nor_606_nl = ~(nor_792_cse | (~ main_stage_v_3));
  assign mux_769_nl = MUX_s_1_2_2(main_stage_v_3, (nor_606_nl), cfg_precision_1_sva_st_70[1]);
  assign mux_1281_nl = MUX_s_1_2_2((mux_769_nl), main_stage_v_3, cfg_precision_1_sva_st_70[0]);
  assign mux_771_cse = (mux_1281_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign nor_609_nl = ~(nor_610_cse | (~ main_stage_v_4));
  assign mux_772_nl = MUX_s_1_2_2(main_stage_v_4, (nor_609_nl), cfg_precision_1_sva_st_71[1]);
  assign mux_773_nl = MUX_s_1_2_2((mux_772_nl), main_stage_v_4, cfg_precision_1_sva_st_71[0]);
  assign mux_774_nl = MUX_s_1_2_2((mux_773_nl), nor_612_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_775_nl = MUX_s_1_2_2((mux_774_nl), mux_771_cse, or_cse);
  assign lut_lookup_if_else_if_and_4_cse = core_wen & (~ and_dcpl_54) & (mux_775_nl);
  assign mux_1187_cse = MUX_s_1_2_2(or_tmp_314, or_1857_cse, or_cse);
  assign nl_lut_lookup_1_IntLog2_32U_acc_1_nl = lut_lookup_1_IntLog2_32U_lshift_itm
      + 31'b1111111111111111111111111111111;
  assign lut_lookup_1_IntLog2_32U_acc_1_nl = nl_lut_lookup_1_IntLog2_32U_acc_1_nl[30:0];
  assign lut_lookup_1_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2
      & (lut_lookup_1_IntLog2_32U_acc_1_nl);
  assign and_649_nl = or_cse & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign lut_lookup_lut_lookup_mux_17_nl = MUX_v_23_2_2((lut_in_data_sva_156[22:0]),
      FpAdd_8U_23U_asn_50_mx0w1, and_649_nl);
  assign IntLog2_32U_mux1h_1_itm = MUX_v_31_2_2(({8'b0 , (lut_lookup_lut_lookup_mux_17_nl)}),
      (lut_lookup_1_IntLog2_32U_and_nl), mux_1187_cse);
  assign and_1142_cse = ((FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp==8'b11111111);
  assign nor_832_cse = ~((~((FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp!=8'b11111111));
  assign nor_434_nl = ~((~ cfg_lut_le_function_1_sva_st_41) | (cfg_precision_1_sva_st_70!=2'b10));
  assign nor_435_nl = ~((~ cfg_lut_le_function_1_sva_st_42) | (cfg_precision_1_sva_st_71!=2'b10));
  assign mux_1188_cse = MUX_s_1_2_2((nor_435_nl), (nor_434_nl), or_cse);
  assign nl_lut_lookup_1_if_else_else_else_else_else_acc_nl = conv_s2u_6_7({1'b1
      , (~ (reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[4:0]))}) + 7'b1011101;
  assign lut_lookup_1_if_else_else_else_else_else_acc_nl = nl_lut_lookup_1_if_else_else_else_else_else_acc_nl[6:0];
  assign nl_lut_lookup_1_if_else_else_else_else_if_acc_nl = ({1'b1 , (reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[4:2])})
      + 4'b1001;
  assign lut_lookup_1_if_else_else_else_else_if_acc_nl = nl_lut_lookup_1_if_else_else_else_else_if_acc_nl[3:0];
  assign nor_432_nl = ~(lut_lookup_1_if_else_else_else_else_acc_itm_32_1 | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_433_nl = ~(cfg_lut_le_function_1_sva_st_42 | lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ or_tmp_314));
  assign mux_1189_nl = MUX_s_1_2_2((nor_433_nl), (nor_432_nl), or_cse);
  assign nor_430_nl = ~((~ lut_lookup_1_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_431_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~(lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      & or_tmp_314)));
  assign mux_1190_nl = MUX_s_1_2_2((nor_431_nl), (nor_430_nl), or_cse);
  assign lut_lookup_else_else_else_else_mux1h_rgt = MUX1HOT_v_9_5_2(lut_lookup_1_else_else_else_else_acc_itm_mx0w0,
      z_out_4, ({1'b0 , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0}),
      ({2'b0 , (lut_lookup_1_if_else_else_else_else_else_acc_nl)}), ({5'b0 , (lut_lookup_1_if_else_else_else_else_if_acc_nl)}),
      {and_dcpl_403 , and_dcpl_405 , mux_1188_cse , (mux_1189_nl) , (mux_1190_nl)});
  assign and_896_cse = (cfg_precision_1_sva_st_70==2'b10);
  assign and_898_cse = (and_896_cse ^ cfg_lut_le_function_1_sva_st_41) & or_cse &
      core_wen;
  assign and_901_cse = (and_896_cse | cfg_lut_le_function_1_sva_st_41) & or_cse &
      core_wen;
  assign and_905_cse = or_cse & core_wen;
  assign and_814_cse = cfg_lut_le_function_1_sva_st_42 & lut_lookup_else_unequal_tmp_18;
  assign and_132_nl = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & lut_lookup_else_else_slc_32_mdf_1_sva_7
      & mux_tmp_704;
  assign mux_1280_nl = MUX_s_1_2_2((and_132_nl), main_stage_v_3, or_1857_cse);
  assign mux_789_cse = (mux_1280_nl) & cfg_lut_le_function_1_sva_st_41;
  assign and_134_cse = cfg_lut_le_function_1_sva_st_42 & main_stage_v_4 & or_tmp_314;
  assign and_653_rgt = or_cse & (~ IsNaN_8U_23U_7_land_1_lpi_1_dfm_7);
  assign nl_lut_lookup_1_else_1_else_else_acc_nl = conv_s2s_8_9(cfg_lut_lo_index_select_1_sva_6)
      + 9'b111011101;
  assign lut_lookup_1_else_1_else_else_acc_nl = nl_lut_lookup_1_else_1_else_else_acc_nl[8:0];
  assign nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl = conv_s2u_7_8(~ (cfg_lut_lo_index_select_1_sva_6[7:1]))
      + 8'b11110101;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl = nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl[7:0];
  assign lut_lookup_else_1_else_else_mux1h_1_itm = MUX_v_9_2_2(({1'b0 , (FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl)}),
      (lut_lookup_1_else_1_else_else_acc_nl), mux_1187_cse);
  assign and_1141_cse = ((FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp==8'b11111111);
  assign mux_805_cse = MUX_s_1_2_2(and_tmp_83, main_stage_v_4, lut_lookup_else_unequal_tmp_18);
  assign nor_588_cse = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (~ FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6)
      | lut_lookup_if_else_else_slc_10_mdf_2_sva_3 | (~(lut_lookup_2_if_else_slc_32_svs_7
      & mux_tmp_704)));
  assign nl_lut_lookup_2_IntLog2_32U_acc_1_nl = lut_lookup_2_IntLog2_32U_lshift_itm
      + 31'b1111111111111111111111111111111;
  assign lut_lookup_2_IntLog2_32U_acc_1_nl = nl_lut_lookup_2_IntLog2_32U_acc_1_nl[30:0];
  assign lut_lookup_2_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1
      & (lut_lookup_2_IntLog2_32U_acc_1_nl);
  assign and_657_nl = or_cse & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign lut_lookup_lut_lookup_mux_nl = MUX_v_23_2_2((lut_in_data_sva_156[54:32]),
      FpAdd_8U_23U_asn_45_mx0w1, and_657_nl);
  assign IntLog2_32U_IntLog2_32U_mux_rgt = MUX_v_31_2_2(({8'b0 , (lut_lookup_lut_lookup_mux_nl)}),
      (lut_lookup_2_IntLog2_32U_and_nl), mux_1187_cse);
  assign and_907_cse = or_cse & core_wen & or_1857_cse;
  assign nl_lut_lookup_2_if_else_else_else_else_else_acc_nl = conv_s2u_6_7({1'b1
      , (~ (reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[4:0]))}) + 7'b1011101;
  assign lut_lookup_2_if_else_else_else_else_else_acc_nl = nl_lut_lookup_2_if_else_else_else_else_else_acc_nl[6:0];
  assign nl_lut_lookup_2_if_else_else_else_else_if_acc_nl = ({1'b1 , (reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[4:2])})
      + 4'b1001;
  assign lut_lookup_2_if_else_else_else_else_if_acc_nl = nl_lut_lookup_2_if_else_else_else_else_if_acc_nl[3:0];
  assign nor_426_nl = ~(lut_lookup_2_if_else_else_else_else_acc_itm_32_1 | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_427_nl = ~(cfg_lut_le_function_1_sva_st_42 | lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ or_tmp_314));
  assign mux_1194_nl = MUX_s_1_2_2((nor_427_nl), (nor_426_nl), or_cse);
  assign nor_424_nl = ~((~ lut_lookup_2_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_425_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~(lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      & or_tmp_314)));
  assign mux_1195_nl = MUX_s_1_2_2((nor_425_nl), (nor_424_nl), or_cse);
  assign lut_lookup_else_else_else_else_mux1h_1_rgt = MUX1HOT_v_9_5_2(lut_lookup_1_else_else_else_else_acc_itm_mx0w0,
      z_out_5, ({1'b0 , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0}),
      ({2'b0 , (lut_lookup_2_if_else_else_else_else_else_acc_nl)}), ({5'b0 , (lut_lookup_2_if_else_else_else_else_if_acc_nl)}),
      {and_dcpl_403 , and_dcpl_405 , mux_1188_cse , (mux_1194_nl) , (mux_1195_nl)});
  assign and_811_cse = cfg_lut_le_function_1_sva_st_42 & lut_lookup_else_unequal_tmp_12;
  assign and_143_nl = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & lut_lookup_else_else_slc_32_mdf_2_sva_7
      & mux_tmp_704;
  assign mux_1279_nl = MUX_s_1_2_2((and_143_nl), main_stage_v_3, or_1857_cse);
  assign mux_845_cse = (mux_1279_nl) & cfg_lut_le_function_1_sva_st_41;
  assign mux_851_cse = MUX_s_1_2_2(and_826_cse, mux_793_cse, cfg_lut_le_function_1_sva_st_41);
  assign mux_852_nl = MUX_s_1_2_2(and_134_cse, main_stage_v_4, and_811_cse);
  assign mux_853_nl = MUX_s_1_2_2((mux_852_nl), mux_851_cse, or_cse);
  assign lut_lookup_else_else_and_5_cse = core_wen & (~ and_dcpl_54) & (mux_853_nl);
  assign and_661_rgt = or_cse & (~ IsNaN_8U_23U_7_land_2_lpi_1_dfm_7);
  assign and_1140_cse = ((FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp==8'b11111111);
  assign nor_564_cse = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (~ FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6)
      | lut_lookup_if_else_else_slc_10_mdf_3_sva_3 | (~(lut_lookup_3_if_else_slc_32_svs_7
      & mux_tmp_704)));
  assign nl_lut_lookup_3_IntLog2_32U_acc_1_nl = lut_lookup_3_IntLog2_32U_lshift_itm
      + 31'b1111111111111111111111111111111;
  assign lut_lookup_3_IntLog2_32U_acc_1_nl = nl_lut_lookup_3_IntLog2_32U_acc_1_nl[30:0];
  assign lut_lookup_3_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1
      & (lut_lookup_3_IntLog2_32U_acc_1_nl);
  assign and_665_nl = or_cse & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign lut_lookup_lut_lookup_mux_3_nl = MUX_v_23_2_2((lut_in_data_sva_156[86:64]),
      FpAdd_8U_23U_asn_40_mx0w1, and_665_nl);
  assign IntLog2_32U_IntLog2_32U_mux_1_rgt = MUX_v_31_2_2(({8'b0 , (lut_lookup_lut_lookup_mux_3_nl)}),
      (lut_lookup_3_IntLog2_32U_and_nl), mux_1187_cse);
  assign nl_lut_lookup_3_if_else_else_else_else_else_acc_nl = conv_s2u_6_7({1'b1
      , (~ (reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[4:0]))}) + 7'b1011101;
  assign lut_lookup_3_if_else_else_else_else_else_acc_nl = nl_lut_lookup_3_if_else_else_else_else_else_acc_nl[6:0];
  assign nl_lut_lookup_3_if_else_else_else_else_if_acc_nl = ({1'b1 , (reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[4:2])})
      + 4'b1001;
  assign lut_lookup_3_if_else_else_else_else_if_acc_nl = nl_lut_lookup_3_if_else_else_else_else_if_acc_nl[3:0];
  assign nor_420_nl = ~(lut_lookup_3_if_else_else_else_else_acc_itm_32_1 | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_421_nl = ~(lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | cfg_lut_le_function_1_sva_st_42 | (~ or_tmp_314));
  assign mux_1199_nl = MUX_s_1_2_2((nor_421_nl), (nor_420_nl), or_cse);
  assign nor_418_nl = ~((~ lut_lookup_3_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_419_nl = ~((~ lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2)
      | cfg_lut_le_function_1_sva_st_42 | (~ or_tmp_314));
  assign mux_1200_nl = MUX_s_1_2_2((nor_419_nl), (nor_418_nl), or_cse);
  assign lut_lookup_else_else_else_else_mux1h_2_rgt = MUX1HOT_v_9_5_2(lut_lookup_1_else_else_else_else_acc_itm_mx0w0,
      z_out_6, ({1'b0 , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0}),
      ({2'b0 , (lut_lookup_3_if_else_else_else_else_else_acc_nl)}), ({5'b0 , (lut_lookup_3_if_else_else_else_else_if_acc_nl)}),
      {and_dcpl_403 , and_dcpl_405 , mux_1188_cse , (mux_1199_nl) , (mux_1200_nl)});
  assign and_153_nl = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & lut_lookup_else_else_slc_32_mdf_3_sva_7
      & mux_tmp_704;
  assign mux_1278_nl = MUX_s_1_2_2((and_153_nl), main_stage_v_3, or_1857_cse);
  assign mux_900_cse = (mux_1278_nl) & cfg_lut_le_function_1_sva_st_41;
  assign and_668_rgt = or_cse & (~ IsNaN_8U_23U_7_land_3_lpi_1_dfm_7);
  assign and_1139_cse = ((FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp==8'b11111111);
  assign mux_917_nl = MUX_s_1_2_2(main_stage_v_4, and_tmp_6, or_cse);
  assign mux_918_nl = MUX_s_1_2_2(and_tmp_83, and_tmp_6, or_cse);
  assign mux_919_nl = MUX_s_1_2_2((mux_918_nl), (mux_917_nl), lut_lookup_else_unequal_tmp_18);
  assign lut_lookup_else_1_and_6_cse = core_wen & (~ and_dcpl_54) & (mux_919_nl);
  assign or_1202_cse = (cfg_precision_1_sva_8!=2'b10);
  assign nl_lut_lookup_4_IntLog2_32U_acc_1_nl = lut_lookup_4_IntLog2_32U_lshift_itm
      + 31'b1111111111111111111111111111111;
  assign lut_lookup_4_IntLog2_32U_acc_1_nl = nl_lut_lookup_4_IntLog2_32U_acc_1_nl[30:0];
  assign lut_lookup_4_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_sva_1
      & (lut_lookup_4_IntLog2_32U_acc_1_nl);
  assign and_672_nl = or_cse & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign lut_lookup_lut_lookup_mux_4_nl = MUX_v_23_2_2((lut_in_data_sva_156[118:96]),
      FpAdd_8U_23U_asn_35_mx0w1, and_672_nl);
  assign IntLog2_32U_IntLog2_32U_mux_2_rgt = MUX_v_31_2_2(({8'b0 , (lut_lookup_lut_lookup_mux_4_nl)}),
      (lut_lookup_4_IntLog2_32U_and_nl), mux_1187_cse);
  assign nl_lut_lookup_4_if_else_else_else_else_else_acc_nl = conv_s2u_6_7({1'b1
      , (~ (reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[4:0]))}) + 7'b1011101;
  assign lut_lookup_4_if_else_else_else_else_else_acc_nl = nl_lut_lookup_4_if_else_else_else_else_else_acc_nl[6:0];
  assign nl_lut_lookup_4_if_else_else_else_else_if_acc_nl = ({1'b1 , (reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[4:2])})
      + 4'b1001;
  assign lut_lookup_4_if_else_else_else_else_if_acc_nl = nl_lut_lookup_4_if_else_else_else_else_if_acc_nl[3:0];
  assign nor_414_nl = ~(lut_lookup_4_if_else_else_else_else_acc_itm_32_1 | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_415_nl = ~(IsNaN_8U_23U_6_land_lpi_1_dfm_6 | (~ or_tmp_314));
  assign mux_1204_nl = MUX_s_1_2_2((nor_415_nl), (nor_414_nl), or_cse);
  assign nor_412_nl = ~((~ lut_lookup_4_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | and_896_cse);
  assign nor_413_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~ IsNaN_8U_23U_6_land_lpi_1_dfm_6));
  assign mux_1205_nl = MUX_s_1_2_2((nor_413_nl), (nor_412_nl), or_cse);
  assign lut_lookup_else_else_else_else_mux1h_3_rgt = MUX1HOT_v_9_5_2(lut_lookup_1_else_else_else_else_acc_itm_mx0w0,
      z_out_7, ({1'b0 , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0}),
      ({2'b0 , (lut_lookup_4_if_else_else_else_else_else_acc_nl)}), ({5'b0 , (lut_lookup_4_if_else_else_else_else_if_acc_nl)}),
      {and_dcpl_403 , and_dcpl_405 , mux_1188_cse , (mux_1204_nl) , (mux_1205_nl)});
  assign nor_526_cse = ~((cfg_precision_1_sva_st_71[1]) | (~ main_stage_v_4));
  assign and_164_nl = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & lut_lookup_else_else_slc_32_mdf_sva_7
      & mux_tmp_704;
  assign mux_1269_nl = MUX_s_1_2_2((and_164_nl), main_stage_v_3, or_1857_cse);
  assign mux_959_cse = (mux_1269_nl) & cfg_lut_le_function_1_sva_st_41;
  assign and_676_rgt = or_cse & (~ IsNaN_8U_23U_7_land_lpi_1_dfm_7);
  assign and_1138_cse = ((FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp==8'b11111111);
  assign lut_lookup_else_and_8_cse = core_wen & lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse
      & mux_tmp_978;
  assign and_679_rgt = (~ or_1857_cse) & or_cse;
  assign and_42_cse = main_stage_v_2 & or_66_cse;
  assign mux_982_cse = MUX_s_1_2_2(and_42_cse, main_stage_v_2, or_66_cse);
  assign and_178_cse = reg_cfg_lut_le_function_1_sva_st_20_cse & mux_982_cse;
  assign and_1179_nl = mux_793_cse & cfg_lut_le_function_1_sva_st_41;
  assign mux_1004_nl = MUX_s_1_2_2((and_1179_nl), and_178_cse, or_cse);
  assign lut_lookup_else_else_and_9_cse = core_wen & (~ and_dcpl_54) & (mux_1004_nl);
  assign mux_1053_nl = MUX_s_1_2_2(and_tmp_6, and_42_cse, or_cse);
  assign lut_lookup_else_1_and_9_cse = core_wen & (~ and_dcpl_54) & (mux_1053_nl);
  assign mux_1056_nl = MUX_s_1_2_2(mux_tmp_704, and_42_cse, or_cse);
  assign lut_lookup_lo_index_0_and_8_cse = core_wen & (~ and_dcpl_54) & (mux_1056_nl);
  assign and_795_cse = (~ IsNaN_8U_23U_3_nor_8_tmp) & (chn_lut_in_rsci_d_mxwt[30:23]==8'b11111111);
  assign and_794_cse = (~ IsNaN_8U_23U_4_nor_tmp) & (cfg_lut_le_start_rsci_d[30:23]==8'b11111111);
  assign and_789_cse = (~ IsNaN_8U_23U_8_nor_2_tmp_1) & (cfg_lut_lo_start_rsci_d[30:23]==8'b11111111);
  assign and_787_cse = (~ IsNaN_8U_23U_3_nor_4_tmp) & (chn_lut_in_rsci_d_mxwt[62:55]==8'b11111111);
  assign and_784_cse = (~ IsNaN_8U_23U_3_nor_10_tmp) & (chn_lut_in_rsci_d_mxwt[94:87]==8'b11111111);
  assign nor_482_cse = ~(IsNaN_8U_23U_8_nor_2_itm_2 | IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2);
  assign nor_478_nl = ~(and_784_cse | (~ chn_lut_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10));
  assign nor_479_nl = ~((~ main_stage_v_1) | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4
      | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign mux_1067_nl = MUX_s_1_2_2((nor_479_nl), (nor_478_nl), or_cse);
  assign IsNaN_8U_23U_8_and_cse = core_wen & (~ and_dcpl_54) & (mux_1067_nl);
  assign and_780_cse = (~ IsNaN_8U_23U_3_nor_6_tmp) & (chn_lut_in_rsci_d_mxwt[126:119]==8'b11111111);
  assign nor_469_cse = ~(IsNaN_8U_23U_8_nor_3_itm_2 | IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2);
  assign nor_465_nl = ~((~ chn_lut_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10)
      | IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0);
  assign nor_466_nl = ~((~ main_stage_v_1) | reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse
      | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign mux_1074_nl = MUX_s_1_2_2((nor_466_nl), (nor_465_nl), or_cse);
  assign IsNaN_8U_23U_8_and_2_cse = core_wen & (~ and_dcpl_54) & (mux_1074_nl);
  assign mux_1106_nl = MUX_s_1_2_2(and_42_cse, mux_tmp_1104, or_cse);
  assign lut_lookup_else_1_and_13_cse = core_wen & (~ and_dcpl_54) & (mux_1106_nl);
  assign mux_1115_nl = MUX_s_1_2_2(mux_tmp_1104, and_tmp_178, or_cse);
  assign lut_lookup_else_1_and_16_cse = core_wen & (~ and_dcpl_54) & (mux_1115_nl);
  assign lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[30:23])
      == (cfg_lut_le_start_rsci_d[30:23]);
  assign lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[30:23])
      == (cfg_lut_lo_start_rsci_d[30:23]);
  assign lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[62:55])
      == (cfg_lut_le_start_rsci_d[30:23]);
  assign lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[62:55])
      == (cfg_lut_lo_start_rsci_d[30:23]);
  assign lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[94:87])
      == (cfg_lut_le_start_rsci_d[30:23]);
  assign lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[94:87])
      == (cfg_lut_lo_start_rsci_d[30:23]);
  assign lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[126:119])
      == (cfg_lut_le_start_rsci_d[30:23]);
  assign lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = (chn_lut_in_rsci_d_mxwt[126:119])
      == (cfg_lut_lo_start_rsci_d[30:23]);
  assign IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_3_nor_8_tmp | (chn_lut_in_rsci_d_mxwt[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_3_nor_6_tmp | (chn_lut_in_rsci_d_mxwt[126:119]!=8'b11111111));
  assign nl_lut_lookup_1_if_else_else_acc_nl = conv_u2u_9_11(signext_9_6({(reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[4:0]))})) - conv_s2u_8_11(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_1_if_else_else_acc_nl = nl_lut_lookup_1_if_else_else_acc_nl[10:0];
  assign lut_lookup_1_if_else_else_acc_itm_10 = readslicef_11_1_10((lut_lookup_1_if_else_else_acc_nl));
  assign FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0 = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[25]));
  assign nl_lut_lookup_1_else_else_else_if_acc_nl = conv_u2u_3_4(IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva[8:6])
      + 4'b1111;
  assign lut_lookup_1_else_else_else_if_acc_nl = nl_lut_lookup_1_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_1_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_1_else_else_else_if_acc_nl));
  assign lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0
      & (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0 = (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[25]));
  assign lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0
      & (FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_lut_lookup_2_if_else_else_acc_nl = conv_u2u_9_11(signext_9_6({(reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[4:0]))})) - conv_s2u_8_11(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_2_if_else_else_acc_nl = nl_lut_lookup_2_if_else_else_acc_nl[10:0];
  assign lut_lookup_2_if_else_else_acc_itm_10 = readslicef_11_1_10((lut_lookup_2_if_else_else_acc_nl));
  assign FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0 = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[25]));
  assign nl_lut_lookup_2_else_else_else_if_acc_nl = conv_u2u_3_4(IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva[8:6])
      + 4'b1111;
  assign lut_lookup_2_else_else_else_if_acc_nl = nl_lut_lookup_2_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_2_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_2_else_else_else_if_acc_nl));
  assign lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0
      & (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0 = (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[25]));
  assign lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0
      & (FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_lut_lookup_3_if_else_else_acc_nl = conv_u2u_9_11(signext_9_6({(reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[4:0]))})) - conv_s2u_8_11(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_3_if_else_else_acc_nl = nl_lut_lookup_3_if_else_else_acc_nl[10:0];
  assign lut_lookup_3_if_else_else_acc_itm_10 = readslicef_11_1_10((lut_lookup_3_if_else_else_acc_nl));
  assign FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0 = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[25]));
  assign nl_lut_lookup_3_else_else_else_if_acc_nl = conv_u2u_3_4(IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva[8:6])
      + 4'b1111;
  assign lut_lookup_3_else_else_else_if_acc_nl = nl_lut_lookup_3_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_3_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_3_else_else_else_if_acc_nl));
  assign lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0
      & (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0 = (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[25]));
  assign lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0
      & (FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_lut_lookup_4_if_else_else_acc_nl = conv_u2u_9_11(signext_9_6({(reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[4:0]))})) - conv_s2u_8_11(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_4_if_else_else_acc_nl = nl_lut_lookup_4_if_else_else_acc_nl[10:0];
  assign lut_lookup_4_if_else_else_acc_itm_10 = readslicef_11_1_10((lut_lookup_4_if_else_else_acc_nl));
  assign FpMantRNE_49U_24U_1_else_carry_sva_mx0w0 = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[25]));
  assign nl_lut_lookup_4_else_else_else_if_acc_nl = conv_u2u_3_4(IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva[8:6])
      + 4'b1111;
  assign lut_lookup_4_else_else_else_if_acc_nl = nl_lut_lookup_4_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_4_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_4_else_else_else_if_acc_nl));
  assign lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_sva_mx0w0
      & (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_2_else_carry_sva_mx0w0 = (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[25]));
  assign lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_sva_mx0w0
      & (FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign nl_lut_lookup_1_if_else_else_else_else_acc_nl = conv_u2s_32_33(signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[4:0]))})) + 33'b111111111111111111111111111011101;
  assign lut_lookup_1_if_else_else_else_else_acc_nl = nl_lut_lookup_1_if_else_else_else_else_acc_nl[32:0];
  assign lut_lookup_1_if_else_else_else_else_acc_itm_32_1 = readslicef_33_1_32((lut_lookup_1_if_else_else_else_else_acc_nl));
  assign lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1 = and_1142_cse | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp
      | FpAdd_8U_23U_1_mux_13_itm_4;
  assign nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0 = conv_s2u_7_8(~
      (cfg_lut_le_index_select_1_sva_6[7:1])) + 8'b11110101;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0 = nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0[7:0];
  assign nl_lut_lookup_1_if_else_else_else_if_acc_nl = conv_u2u_3_4({reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
      , reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm})
      + 4'b1111;
  assign lut_lookup_1_if_else_else_else_if_acc_nl = nl_lut_lookup_1_if_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_1_if_else_else_else_if_acc_itm_3 = readslicef_4_1_3((lut_lookup_1_if_else_else_else_if_acc_nl));
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp = ~((FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp!=8'b00000000));
  assign nl_lut_lookup_2_if_else_else_else_else_acc_nl = conv_u2s_32_33(signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[4:0]))})) + 33'b111111111111111111111111111011101;
  assign lut_lookup_2_if_else_else_else_else_acc_nl = nl_lut_lookup_2_if_else_else_else_else_acc_nl[32:0];
  assign lut_lookup_2_if_else_else_else_else_acc_itm_32_1 = readslicef_33_1_32((lut_lookup_2_if_else_else_else_else_acc_nl));
  assign lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1 = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp | FpAdd_8U_23U_1_mux_29_itm_4;
  assign nl_lut_lookup_2_if_else_else_else_if_acc_nl = conv_u2u_3_4({reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
      , reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm})
      + 4'b1111;
  assign lut_lookup_2_if_else_else_else_if_acc_nl = nl_lut_lookup_2_if_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_2_if_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_2_if_else_else_else_if_acc_nl));
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp = ~((FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp!=8'b00000000));
  assign lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0 = and_1140_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp
      | FpAdd_8U_23U_2_mux_29_itm_3;
  assign nl_lut_lookup_3_if_else_else_else_else_acc_nl = conv_u2s_32_33(signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[4:0]))})) + 33'b111111111111111111111111111011101;
  assign lut_lookup_3_if_else_else_else_else_acc_nl = nl_lut_lookup_3_if_else_else_else_else_acc_nl[32:0];
  assign lut_lookup_3_if_else_else_else_else_acc_itm_32_1 = readslicef_33_1_32((lut_lookup_3_if_else_else_else_else_acc_nl));
  assign lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1 = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp | FpAdd_8U_23U_1_mux_45_itm_4;
  assign nl_lut_lookup_3_if_else_else_else_if_acc_nl = conv_u2u_3_4({reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
      , reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm})
      + 4'b1111;
  assign lut_lookup_3_if_else_else_else_if_acc_nl = nl_lut_lookup_3_if_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_3_if_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_3_if_else_else_else_if_acc_nl));
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp = ~((FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp!=8'b00000000));
  assign lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0 = and_1139_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp
      | FpAdd_8U_23U_2_mux_45_itm_3;
  assign nl_lut_lookup_4_if_else_else_else_else_acc_nl = conv_u2s_32_33(signext_32_6({(reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[4:0]))})) + 33'b111111111111111111111111111011101;
  assign lut_lookup_4_if_else_else_else_else_acc_nl = nl_lut_lookup_4_if_else_else_else_else_acc_nl[32:0];
  assign lut_lookup_4_if_else_else_else_else_acc_itm_32_1 = readslicef_33_1_32((lut_lookup_4_if_else_else_else_else_acc_nl));
  assign lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1 = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp
      | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp | FpAdd_8U_23U_1_mux_61_itm_4;
  assign nl_lut_lookup_4_if_else_else_else_if_acc_nl = conv_u2u_3_4({reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
      , reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm})
      + 4'b1111;
  assign lut_lookup_4_if_else_else_else_if_acc_nl = nl_lut_lookup_4_if_else_else_else_if_acc_nl[3:0];
  assign lut_lookup_4_if_else_else_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_4_if_else_else_else_if_acc_nl));
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp = ~((FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp!=8'b00000000));
  assign lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0 = and_1138_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp
      | FpAdd_8U_23U_2_mux_61_itm_3;
  assign lut_lookup_if_unequal_tmp_1_mx0w0 = ~((cfg_precision_1_sva_8==2'b10));
  assign lut_lookup_if_else_lut_lookup_if_else_or_3_cse = lut_lookup_if_else_else_slc_10_mdf_sva_4
      | (~ lut_lookup_4_if_else_slc_32_svs_8);
  assign lut_lookup_if_if_lut_lookup_if_if_or_3_nl = lut_lookup_4_if_if_else_acc_itm_9_1
      | lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  assign lut_lookup_if_mux_123_mx0w1 = MUX_s_1_2_2((lut_lookup_if_if_lut_lookup_if_if_or_3_nl),
      lut_lookup_if_else_lut_lookup_if_else_or_3_cse, lut_lookup_if_unequal_tmp_1_mx0w0);
  assign lut_lookup_if_else_lut_lookup_if_else_or_2_cse = lut_lookup_if_else_else_slc_10_mdf_3_sva_4
      | (~ lut_lookup_3_if_else_slc_32_svs_8);
  assign lut_lookup_if_if_lut_lookup_if_if_or_2_nl = lut_lookup_3_if_if_else_acc_itm_9_1
      | lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  assign lut_lookup_if_mux_82_mx0w1 = MUX_s_1_2_2((lut_lookup_if_if_lut_lookup_if_if_or_2_nl),
      lut_lookup_if_else_lut_lookup_if_else_or_2_cse, lut_lookup_if_unequal_tmp_1_mx0w0);
  assign lut_lookup_if_else_lut_lookup_if_else_or_1_cse = lut_lookup_if_else_else_slc_10_mdf_2_sva_4
      | (~ lut_lookup_2_if_else_slc_32_svs_8);
  assign lut_lookup_if_if_lut_lookup_if_if_or_1_nl = lut_lookup_2_if_if_else_acc_itm_9_1
      | lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  assign lut_lookup_if_mux_41_mx0w1 = MUX_s_1_2_2((lut_lookup_if_if_lut_lookup_if_if_or_1_nl),
      lut_lookup_if_else_lut_lookup_if_else_or_1_cse, lut_lookup_if_unequal_tmp_1_mx0w0);
  assign lut_lookup_if_else_lut_lookup_if_else_or_cse = lut_lookup_if_else_else_slc_10_mdf_1_sva_4
      | (~ lut_lookup_1_if_else_slc_32_svs_8);
  assign lut_lookup_if_if_lut_lookup_if_if_or_nl = lut_lookup_1_if_if_else_acc_itm_9_1
      | lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  assign lut_lookup_if_mux_mx0w1 = MUX_s_1_2_2((lut_lookup_if_if_lut_lookup_if_if_or_nl),
      lut_lookup_if_else_lut_lookup_if_else_or_cse, lut_lookup_if_unequal_tmp_1_mx0w0);
  assign lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = (cfg_lut_le_start_rsci_d[30:0]!=31'b0000000000000000000000000000000);
  assign lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = (chn_lut_in_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000);
  assign nl_lut_lookup_1_else_1_acc_nl = conv_s2u_32_33(cfg_lut_lo_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[31:0]);
  assign lut_lookup_1_else_1_acc_nl = nl_lut_lookup_1_else_1_acc_nl[32:0];
  assign lut_lookup_1_else_1_acc_itm_32 = readslicef_33_1_32((lut_lookup_1_else_1_acc_nl));
  assign lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = (chn_lut_in_rsci_d_mxwt[62:32]!=31'b0000000000000000000000000000000);
  assign nl_lut_lookup_2_else_1_acc_nl = conv_s2u_32_33(cfg_lut_lo_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[63:32]);
  assign lut_lookup_2_else_1_acc_nl = nl_lut_lookup_2_else_1_acc_nl[32:0];
  assign lut_lookup_2_else_1_acc_itm_32 = readslicef_33_1_32((lut_lookup_2_else_1_acc_nl));
  assign lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = (chn_lut_in_rsci_d_mxwt[94:64]!=31'b0000000000000000000000000000000);
  assign nl_lut_lookup_3_else_1_acc_nl = conv_s2u_32_33(cfg_lut_lo_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[95:64]);
  assign lut_lookup_3_else_1_acc_nl = nl_lut_lookup_3_else_1_acc_nl[32:0];
  assign lut_lookup_3_else_1_acc_itm_32 = readslicef_33_1_32((lut_lookup_3_else_1_acc_nl));
  assign lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = (chn_lut_in_rsci_d_mxwt[126:96]!=31'b0000000000000000000000000000000);
  assign nl_lut_lookup_4_else_1_acc_nl = conv_s2u_32_33(cfg_lut_lo_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[127:96]);
  assign lut_lookup_4_else_1_acc_nl = nl_lut_lookup_4_else_1_acc_nl[32:0];
  assign lut_lookup_4_else_1_acc_itm_32 = readslicef_33_1_32((lut_lookup_4_else_1_acc_nl));
  assign IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_4_nor_3_itm_2 | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2);
  assign IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_4_nor_itm_2 | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2);
  assign nl_lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0 = (lut_in_data_sva_154[31:0])
      - cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0 = nl_lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0[31:0];
  assign nl_lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0 = (lut_in_data_sva_154[63:32])
      - cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0 = nl_lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0[31:0];
  assign nl_lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0 = (lut_in_data_sva_154[95:64])
      - cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0 = nl_lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0[31:0];
  assign nl_lut_lookup_if_else_else_le_data_sub_sva_mx0w0 = (lut_in_data_sva_154[127:96])
      - cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_sva_mx0w0 = nl_lut_lookup_if_else_else_le_data_sub_sva_mx0w0[31:0];
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp = ((FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_o_expo_lpi_1_dfm_7==8'b11111111);
  assign lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3 = (~((~((FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_o_expo_lpi_1_dfm_7!=8'b11111111))) | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp
      | FpAdd_8U_23U_1_mux_61_itm_4;
  assign lut_lookup_unequal_tmp_mx0w0 = ~((cfg_precision_1_sva_st_70==2'b10));
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp = ((FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7==8'b11111111);
  assign lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3 = (~((~((FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7!=8'b11111111))) | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp
      | FpAdd_8U_23U_1_mux_45_itm_4;
  assign lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3 = (~((~((FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7!=8'b11111111))) | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp
      | FpAdd_8U_23U_1_mux_29_itm_4;
  assign lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3 = nor_832_cse | IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp
      | FpAdd_8U_23U_1_mux_13_itm_4;
  assign nl_lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_1_else_carry_1_sva_2);
  assign lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl = nl_lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl = MUX_v_23_2_2((lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_asn_50_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl),
      (cfg_lut_le_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_1_land_1_lpi_1_dfm_8);
  assign nl_lut_lookup_1_else_else_else_else_acc_itm_mx0w0 = conv_s2s_8_9(cfg_lut_le_index_select_1_sva_6)
      + 9'b111011101;
  assign lut_lookup_1_else_else_else_else_acc_itm_mx0w0 = nl_lut_lookup_1_else_else_else_else_acc_itm_mx0w0[8:0];
  assign nl_lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_2_else_carry_1_sva_2);
  assign lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl = nl_lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl[22:0];
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_4_nl = MUX_v_23_2_2((lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_2_asn_50_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_4_nl),
      (cfg_lut_lo_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_8_land_2_lpi_1_dfm_7);
  assign nl_lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_1_else_carry_2_sva_2);
  assign lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl = nl_lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl = MUX_v_23_2_2((lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_asn_45_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl),
      (cfg_lut_le_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_1_land_2_lpi_1_dfm_8);
  assign nl_lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_2_else_carry_2_sva_2);
  assign lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl = nl_lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl[22:0];
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_5_nl = MUX_v_23_2_2((lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_2_asn_45_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_5_nl),
      (cfg_lut_lo_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_8_land_2_lpi_1_dfm_7);
  assign nl_lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_1_else_carry_3_sva_2);
  assign lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl = nl_lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl = MUX_v_23_2_2((lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_asn_40_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl),
      (cfg_lut_le_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_1_land_3_lpi_1_dfm_8);
  assign nl_lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_2_else_carry_3_sva_2);
  assign lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl = nl_lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl[22:0];
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_6_nl = MUX_v_23_2_2((lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_2_asn_40_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_6_nl),
      (cfg_lut_lo_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_8_land_3_lpi_1_dfm_5);
  assign nl_lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_1_else_carry_sva_2);
  assign lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl = nl_lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl = MUX_v_23_2_2((lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_asn_35_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl),
      (cfg_lut_le_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_1_land_lpi_1_dfm_8);
  assign nl_lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
      + conv_u2u_1_23(FpMantRNE_49U_24U_2_else_carry_sva_2);
  assign lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl = nl_lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl[22:0];
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_7_nl = MUX_v_23_2_2((lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_2_asn_35_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_7_nl),
      (cfg_lut_lo_start_1_sva_3_30_0_1[22:0]), IsNaN_8U_23U_8_land_lpi_1_dfm_5);
  assign IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_4_nor_tmp | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0);
  assign IsNaN_8U_23U_4_nor_tmp = ~((cfg_lut_le_start_rsci_d[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0 = ~((cfg_lut_le_start_rsci_d[30:23]==8'b11111111));
  assign IsNaN_8U_23U_8_nor_2_tmp_1 = ~((cfg_lut_lo_start_rsci_d[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0 = ~((cfg_lut_lo_start_rsci_d[30:23]==8'b11111111));
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_nl = ({1'b1 , (cfg_lut_lo_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[30:23])) + 9'b1;
  assign FpAdd_8U_23U_2_is_a_greater_acc_nl = nl_FpAdd_8U_23U_2_is_a_greater_acc_nl[8:0];
  assign FpAdd_8U_23U_2_is_a_greater_acc_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_2_is_a_greater_acc_nl));
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_1_nl = ({1'b1 , (cfg_lut_lo_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[62:55])) + 9'b1;
  assign FpAdd_8U_23U_2_is_a_greater_acc_1_nl = nl_FpAdd_8U_23U_2_is_a_greater_acc_1_nl[8:0];
  assign FpAdd_8U_23U_2_is_a_greater_acc_1_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_2_is_a_greater_acc_1_nl));
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_2_nl = ({1'b1 , (cfg_lut_lo_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[94:87])) + 9'b1;
  assign FpAdd_8U_23U_2_is_a_greater_acc_2_nl = nl_FpAdd_8U_23U_2_is_a_greater_acc_2_nl[8:0];
  assign FpAdd_8U_23U_2_is_a_greater_acc_2_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_2_is_a_greater_acc_2_nl));
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_3_nl = ({1'b1 , (cfg_lut_lo_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[126:119])) + 9'b1;
  assign FpAdd_8U_23U_2_is_a_greater_acc_3_nl = nl_FpAdd_8U_23U_2_is_a_greater_acc_3_nl[8:0];
  assign FpAdd_8U_23U_2_is_a_greater_acc_3_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_2_is_a_greater_acc_3_nl));
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5[7:1])})
      + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0];
  assign lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl));
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5[7:1])})
      + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0];
  assign lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl));
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5[7:1])})
      + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0];
  assign lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl));
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_qr_lpi_1_dfm_5[7:1])})
      + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0];
  assign lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6
      | (~ lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl), reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse);
  assign FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_asn_50_mx0w1,
      (lut_in_data_sva_156[22:0]), IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign nl_lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl = ({reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm}) + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_59_nl = (~(FpAdd_8U_23U_1_and_tmp | FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_and_61_nl = FpAdd_8U_23U_1_and_tmp & (~ FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_1_and_35_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_and_35_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp = MUX1HOT_v_8_5_2(({reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm}), (lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl),
      8'b11111110, (cfg_lut_le_start_1_sva_3_30_0_1[30:23]), (lut_in_data_sva_156[30:23]),
      {(FpAdd_8U_23U_and_59_nl) , (FpAdd_8U_23U_and_61_nl) , (FpAdd_8U_23U_1_and_35_nl)
      , (FpAdd_8U_23U_and_35_nl) , IsNaN_8U_23U_3_land_1_lpi_1_dfm_6});
  assign FpAdd_8U_23U_1_and_tmp = lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1
      & reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12[7:1])})
      + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0];
  assign lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_4_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5
      | (~ lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5,
      (FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_4_nl), lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_2_asn_50_mx0w1,
      (lut_in_data_sva_156[22:0]), IsNaN_8U_23U_7_land_1_lpi_1_dfm_7);
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12
      + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_2_and_nl = (~(FpAdd_8U_23U_2_and_tmp | FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  assign FpAdd_8U_23U_2_and_6_nl = FpAdd_8U_23U_2_and_tmp & (~ FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  assign FpAdd_8U_23U_2_and_28_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  assign FpAdd_8U_23U_2_and_9_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 & (~ IsNaN_8U_23U_7_land_1_lpi_1_dfm_7);
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp = MUX1HOT_v_8_5_2(FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12,
      (lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl), 8'b11111110, (cfg_lut_lo_start_1_sva_3_30_0_1[30:23]),
      (lut_in_data_sva_156[30:23]), {(FpAdd_8U_23U_2_and_nl) , (FpAdd_8U_23U_2_and_6_nl)
      , (FpAdd_8U_23U_2_and_28_nl) , (FpAdd_8U_23U_2_and_9_nl) , IsNaN_8U_23U_7_land_1_lpi_1_dfm_7});
  assign FpAdd_8U_23U_2_and_tmp = lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1
      & lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c = ~(IsNaN_8U_23U_8_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_7_land_1_lpi_1_dfm_7);
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6
      | (~ lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl), reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse);
  assign FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_asn_45_mx0w1,
      (lut_in_data_sva_156[54:32]), IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign nl_lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl = ({reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm}) + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_63_nl = (~(FpAdd_8U_23U_1_and_1_tmp | FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_and_65_nl = FpAdd_8U_23U_1_and_1_tmp & (~ FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_1_and_37_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_and_37_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7 = MUX1HOT_v_8_5_2(({reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm}), (lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl),
      8'b11111110, (cfg_lut_le_start_1_sva_3_30_0_1[30:23]), (lut_in_data_sva_156[62:55]),
      {(FpAdd_8U_23U_and_63_nl) , (FpAdd_8U_23U_and_65_nl) , (FpAdd_8U_23U_1_and_37_nl)
      , (FpAdd_8U_23U_and_37_nl) , IsNaN_8U_23U_3_land_2_lpi_1_dfm_7});
  assign FpAdd_8U_23U_1_and_1_tmp = lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1
      & reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp = ((FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0!=23'b00000000000000000000000))
      & (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7==8'b11111111);
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12[7:1])})
      + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0];
  assign lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_5_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5
      | (~ lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5,
      (FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_5_nl), lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_2_asn_45_mx0w1,
      (lut_in_data_sva_156[54:32]), IsNaN_8U_23U_7_land_2_lpi_1_dfm_7);
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12
      + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_2_and_29_nl = (~(FpAdd_8U_23U_2_and_1_tmp | FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  assign FpAdd_8U_23U_2_and_13_nl = FpAdd_8U_23U_2_and_1_tmp & (~ FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  assign FpAdd_8U_23U_2_and_30_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  assign FpAdd_8U_23U_2_and_15_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 & (~ IsNaN_8U_23U_7_land_2_lpi_1_dfm_7);
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp = MUX1HOT_v_8_5_2(FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12,
      (lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl), 8'b11111110, (cfg_lut_lo_start_1_sva_3_30_0_1[30:23]),
      (lut_in_data_sva_156[62:55]), {(FpAdd_8U_23U_2_and_29_nl) , (FpAdd_8U_23U_2_and_13_nl)
      , (FpAdd_8U_23U_2_and_30_nl) , (FpAdd_8U_23U_2_and_15_nl) , IsNaN_8U_23U_7_land_2_lpi_1_dfm_7});
  assign FpAdd_8U_23U_2_and_1_tmp = lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1
      & lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c = ~(IsNaN_8U_23U_8_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_7_land_2_lpi_1_dfm_7);
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6
      | (~ lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl), reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse);
  assign FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_asn_40_mx0w1,
      (lut_in_data_sva_156[86:64]), IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign nl_lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl = ({reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm}) + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_67_nl = (~(FpAdd_8U_23U_1_and_2_tmp | FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_and_69_nl = FpAdd_8U_23U_1_and_2_tmp & (~ FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_1_and_39_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_and_39_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7 = MUX1HOT_v_8_5_2(({reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm}), (lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl),
      8'b11111110, (cfg_lut_le_start_1_sva_3_30_0_1[30:23]), (lut_in_data_sva_156[94:87]),
      {(FpAdd_8U_23U_and_67_nl) , (FpAdd_8U_23U_and_69_nl) , (FpAdd_8U_23U_1_and_39_nl)
      , (FpAdd_8U_23U_and_39_nl) , IsNaN_8U_23U_3_land_3_lpi_1_dfm_7});
  assign FpAdd_8U_23U_1_and_2_tmp = lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1
      & reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12[7:1])})
      + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0];
  assign lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_6_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5
      | (~ lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5,
      (FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_6_nl), lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_2_asn_40_mx0w1,
      (lut_in_data_sva_156[86:64]), IsNaN_8U_23U_7_land_3_lpi_1_dfm_7);
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12
      + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_2_and_31_nl = (~(FpAdd_8U_23U_2_and_2_tmp | FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  assign FpAdd_8U_23U_2_and_19_nl = FpAdd_8U_23U_2_and_2_tmp & (~ FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  assign FpAdd_8U_23U_2_and_32_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  assign FpAdd_8U_23U_2_and_21_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 & (~ IsNaN_8U_23U_7_land_3_lpi_1_dfm_7);
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp = MUX1HOT_v_8_5_2(FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12,
      (lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl), 8'b11111110, (cfg_lut_lo_start_1_sva_3_30_0_1[30:23]),
      (lut_in_data_sva_156[94:87]), {(FpAdd_8U_23U_2_and_31_nl) , (FpAdd_8U_23U_2_and_19_nl)
      , (FpAdd_8U_23U_2_and_32_nl) , (FpAdd_8U_23U_2_and_21_nl) , IsNaN_8U_23U_7_land_3_lpi_1_dfm_7});
  assign FpAdd_8U_23U_2_and_2_tmp = lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1
      & lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c = ~(IsNaN_8U_23U_8_land_3_lpi_1_dfm_5
      | IsNaN_8U_23U_7_land_3_lpi_1_dfm_7);
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6
      | (~ lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl), reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse);
  assign FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_asn_35_mx0w1,
      (lut_in_data_sva_156[118:96]), IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign nl_lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl = ({reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm}) + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_71_nl = (~(FpAdd_8U_23U_1_and_3_tmp | FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_and_73_nl = FpAdd_8U_23U_1_and_3_tmp & (~ FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_1_and_41_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_and_41_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_8 & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_7 = MUX1HOT_v_8_5_2(({reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm
      , reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm}), (lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl),
      8'b11111110, (cfg_lut_le_start_1_sva_3_30_0_1[30:23]), (lut_in_data_sva_156[126:119]),
      {(FpAdd_8U_23U_and_71_nl) , (FpAdd_8U_23U_and_73_nl) , (FpAdd_8U_23U_1_and_41_nl)
      , (FpAdd_8U_23U_and_41_nl) , IsNaN_8U_23U_3_land_lpi_1_dfm_6});
  assign FpAdd_8U_23U_1_and_3_tmp = lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1
      & reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12[7:1])})
      + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0];
  assign lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_7_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5
      | (~ lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5,
      (FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_7_nl), lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0 = MUX_v_23_2_2(FpAdd_8U_23U_2_asn_35_mx0w1,
      (lut_in_data_sva_156[118:96]), IsNaN_8U_23U_7_land_lpi_1_dfm_7);
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12
      + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_2_and_33_nl = (~(FpAdd_8U_23U_2_and_3_tmp | FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  assign FpAdd_8U_23U_2_and_25_nl = FpAdd_8U_23U_2_and_3_tmp & (~ FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  assign FpAdd_8U_23U_2_and_34_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  assign FpAdd_8U_23U_2_and_27_nl = IsNaN_8U_23U_8_land_lpi_1_dfm_5 & (~ IsNaN_8U_23U_7_land_lpi_1_dfm_7);
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp = MUX1HOT_v_8_5_2(FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12,
      (lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl), 8'b11111110, (cfg_lut_lo_start_1_sva_3_30_0_1[30:23]),
      (lut_in_data_sva_156[126:119]), {(FpAdd_8U_23U_2_and_33_nl) , (FpAdd_8U_23U_2_and_25_nl)
      , (FpAdd_8U_23U_2_and_34_nl) , (FpAdd_8U_23U_2_and_27_nl) , IsNaN_8U_23U_7_land_lpi_1_dfm_7});
  assign FpAdd_8U_23U_2_and_3_tmp = lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1
      & lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c = ~(IsNaN_8U_23U_8_land_lpi_1_dfm_5
      | IsNaN_8U_23U_7_land_lpi_1_dfm_7);
  assign nl_lut_lookup_1_if_if_else_acc_nl = conv_s2u_9_10({reg_lut_lookup_1_else_else_else_else_acc_reg
      , reg_lut_lookup_1_else_else_else_else_acc_1_reg , reg_lut_lookup_1_else_else_else_else_acc_2_reg
      , reg_lut_lookup_1_else_else_else_else_acc_3_reg}) - conv_s2u_8_10(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_1_if_if_else_acc_nl = nl_lut_lookup_1_if_if_else_acc_nl[9:0];
  assign lut_lookup_1_if_if_else_acc_itm_9_1 = readslicef_10_1_9((lut_lookup_1_if_if_else_acc_nl));
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_1_else_else_else_else_acc_1_reg
      , reg_lut_lookup_1_else_else_else_else_acc_2_reg , reg_lut_lookup_1_else_else_else_else_acc_3_reg
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2);
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_1_else_1_else_else_acc_1_itm
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2);
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_2_if_if_else_acc_nl = conv_s2u_9_10({reg_lut_lookup_2_else_else_else_else_acc_reg
      , reg_lut_lookup_2_else_else_else_else_acc_1_reg , reg_lut_lookup_2_else_else_else_else_acc_2_reg
      , reg_lut_lookup_2_else_else_else_else_acc_3_reg}) - conv_s2u_8_10(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_2_if_if_else_acc_nl = nl_lut_lookup_2_if_if_else_acc_nl[9:0];
  assign lut_lookup_2_if_if_else_acc_itm_9_1 = readslicef_10_1_9((lut_lookup_2_if_if_else_acc_nl));
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_2_else_else_else_else_acc_1_reg
      , reg_lut_lookup_2_else_else_else_else_acc_2_reg , reg_lut_lookup_2_else_else_else_else_acc_3_reg
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2);
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_2_else_1_else_else_acc_1_itm
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2);
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_3_if_if_else_acc_nl = conv_s2u_9_10({reg_lut_lookup_3_else_else_else_else_acc_reg
      , reg_lut_lookup_3_else_else_else_else_acc_1_reg , reg_lut_lookup_3_else_else_else_else_acc_2_reg
      , reg_lut_lookup_3_else_else_else_else_acc_3_reg}) - conv_s2u_8_10(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_3_if_if_else_acc_nl = nl_lut_lookup_3_if_if_else_acc_nl[9:0];
  assign lut_lookup_3_if_if_else_acc_itm_9_1 = readslicef_10_1_9((lut_lookup_3_if_if_else_acc_nl));
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_3_else_else_else_else_acc_1_reg
      , reg_lut_lookup_3_else_else_else_else_acc_2_reg , reg_lut_lookup_3_else_else_else_else_acc_3_reg
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2);
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_3_else_1_else_else_acc_1_itm
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2);
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_4_if_if_else_acc_nl = conv_s2u_9_10({reg_lut_lookup_4_else_else_else_else_acc_reg
      , reg_lut_lookup_4_else_else_else_else_acc_1_reg , reg_lut_lookup_4_else_else_else_else_acc_2_reg
      , reg_lut_lookup_4_else_else_else_else_acc_3_reg}) - conv_s2u_8_10(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_4_if_if_else_acc_nl = nl_lut_lookup_4_if_if_else_acc_nl[9:0];
  assign lut_lookup_4_if_if_else_acc_itm_9_1 = readslicef_10_1_9((lut_lookup_4_if_if_else_acc_nl));
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_4_else_else_else_else_acc_1_reg
      , reg_lut_lookup_4_else_else_else_else_acc_2_reg , reg_lut_lookup_4_else_else_else_else_acc_3_reg
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2);
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = conv_s2s_9_10({reg_lut_lookup_4_else_1_else_else_acc_1_itm
      , FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1}) + conv_s2s_8_10(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2);
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0];
  assign nl_lut_lookup_1_else_if_else_if_acc_nl = conv_u2u_3_4(lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1[8:6])
      + 4'b1111;
  assign lut_lookup_1_else_if_else_if_acc_nl = nl_lut_lookup_1_else_if_else_if_acc_nl[3:0];
  assign lut_lookup_1_else_if_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_1_else_if_else_if_acc_nl));
  assign lut_lookup_lo_miss_1_sva = lut_lookup_lo_uflow_1_lpi_1_dfm_4 | lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse
      = lut_lookup_lo_miss_1_sva & lut_lookup_le_miss_1_sva;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_nl = ~(lut_lookup_1_else_if_else_if_acc_itm_3_1
      | lut_lookup_else_if_lor_5_lpi_1_dfm_6);
  assign lut_lookup_else_mux_172_nl = MUX_s_1_2_2((lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_nl),
      lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2, lut_lookup_unequal_tmp_13);
  assign lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0 = MUX_s_1_2_2(lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2,
      (lut_lookup_else_mux_172_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_if_1_lut_lookup_if_1_and_11_nl = (lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[8])
      & (~ lut_lookup_if_1_lor_5_lpi_1_dfm_5);
  assign lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2((lut_lookup_if_1_lut_lookup_if_1_and_11_nl),
      lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2, lut_lookup_unequal_tmp_13);
  assign lut_lookup_le_miss_1_sva = lut_lookup_le_uflow_1_lpi_1_dfm_6 | lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6 = MUX_v_2_2_2((lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1[7:6]),
      (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13[7:6]), lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_mux_2_cse_mx0 = MUX_s_1_2_2(lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse = (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~(lut_lookup_le_miss_1_sva
      | lut_lookup_lo_miss_1_sva);
  assign lut_lookup_le_fraction_1_lpi_1_dfm_9 = lut_lookup_else_if_else_le_fra_1_sva_4
      & ({{34{lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2}},
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_6_land_1_lpi_1_dfm_7)) & ({{34{lut_lookup_1_else_if_else_if_acc_itm_3_1}},
      lut_lookup_1_else_if_else_if_acc_itm_3_1}) & (signext_35_1(~ lut_lookup_else_if_lor_5_lpi_1_dfm_6));
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = ({1'b1 ,
      (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2[8:0]),
      9'b111111111, (readslicef_248_1_247((lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl)))));
  assign lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_nl),
      9'b111111111, IsNaN_8U_23U_6_land_1_lpi_1_dfm_7));
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = ({1'b1
      , (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0];
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = readslicef_248_1_247((lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl));
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2[8:0]),
      9'b111111111, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1));
  assign lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_nl),
      9'b111111111, IsNaN_8U_23U_10_land_1_lpi_1_dfm_6));
  assign lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1 = (lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[7:0])
      & (signext_8_1(~ (lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[8]))) & (signext_8_1(~
      lut_lookup_if_1_lor_5_lpi_1_dfm_5));
  assign lut_lookup_lo_fraction_1_lpi_1_dfm_1 = lut_lookup_if_1_else_lo_fra_1_sva_4
      & ({{34{lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2}},
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_10_land_1_lpi_1_dfm_6)) & (signext_35_1(~ (lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[8])))
      & (signext_35_1(~ lut_lookup_if_1_lor_5_lpi_1_dfm_5));
  assign lut_lookup_1_else_2_and_svs = lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0
      & lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0;
  assign nl_lut_lookup_2_else_if_else_if_acc_nl = conv_u2u_3_4(lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1[8:6])
      + 4'b1111;
  assign lut_lookup_2_else_if_else_if_acc_nl = nl_lut_lookup_2_else_if_else_if_acc_nl[3:0];
  assign lut_lookup_2_else_if_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_2_else_if_else_if_acc_nl));
  assign lut_lookup_lo_miss_2_sva = lut_lookup_lo_uflow_2_lpi_1_dfm_4 | lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_2_sva = lut_lookup_le_uflow_2_lpi_1_dfm_6 | lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse
      = lut_lookup_lo_miss_2_sva & lut_lookup_le_miss_2_sva;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_1_nl = ~(lut_lookup_2_else_if_else_if_acc_itm_3_1
      | lut_lookup_else_if_lor_6_lpi_1_dfm_6);
  assign lut_lookup_else_mux_174_nl = MUX_s_1_2_2((lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_1_nl),
      lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2, lut_lookup_else_unequal_tmp_13);
  assign lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0 = MUX_s_1_2_2(lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2,
      (lut_lookup_else_mux_174_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_if_1_lut_lookup_if_1_and_12_nl = (lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[8])
      & (~ lut_lookup_if_1_lor_6_lpi_1_dfm_5);
  assign lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2((lut_lookup_if_1_lut_lookup_if_1_and_12_nl),
      lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2, lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6 = MUX_v_2_2_2((lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1[7:6]),
      (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13[7:6]), lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse = (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_mux_7_cse_mx0 = MUX_s_1_2_2(lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~(lut_lookup_le_miss_2_sva
      | lut_lookup_lo_miss_2_sva);
  assign lut_lookup_le_fraction_2_lpi_1_dfm_9 = lut_lookup_else_if_else_le_fra_2_sva_4
      & ({{34{lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2}},
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_6_land_2_lpi_1_dfm_7)) & ({{34{lut_lookup_2_else_if_else_if_acc_itm_3_1}},
      lut_lookup_2_else_if_else_if_acc_itm_3_1}) & (signext_35_1(~ lut_lookup_else_if_lor_6_lpi_1_dfm_6));
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = ({1'b1 ,
      (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_1_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2[8:0]),
      9'b111111111, (readslicef_248_1_247((lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl)))));
  assign lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_1_nl),
      9'b111111111, IsNaN_8U_23U_6_land_2_lpi_1_dfm_7));
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = ({1'b1
      , (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0];
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = readslicef_248_1_247((lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl));
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_1_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2[8:0]),
      9'b111111111, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1));
  assign lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_1_nl),
      9'b111111111, IsNaN_8U_23U_10_land_2_lpi_1_dfm_6));
  assign lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1 = (lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[7:0])
      & (signext_8_1(~ (lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[8]))) & (signext_8_1(~
      lut_lookup_if_1_lor_6_lpi_1_dfm_5));
  assign lut_lookup_lo_fraction_2_lpi_1_dfm_1 = lut_lookup_if_1_else_lo_fra_2_sva_4
      & ({{34{lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2}},
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_10_land_2_lpi_1_dfm_6)) & (signext_35_1(~ (lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[8])))
      & (signext_35_1(~ lut_lookup_if_1_lor_6_lpi_1_dfm_5));
  assign lut_lookup_2_else_2_and_svs = lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0
      & lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0;
  assign nl_lut_lookup_3_else_if_else_if_acc_nl = conv_u2u_3_4(lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1[8:6])
      + 4'b1111;
  assign lut_lookup_3_else_if_else_if_acc_nl = nl_lut_lookup_3_else_if_else_if_acc_nl[3:0];
  assign lut_lookup_3_else_if_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_3_else_if_else_if_acc_nl));
  assign lut_lookup_lo_miss_3_sva = lut_lookup_lo_uflow_3_lpi_1_dfm_4 | lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_3_sva = lut_lookup_le_uflow_3_lpi_1_dfm_6 | lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse
      = lut_lookup_lo_miss_3_sva & lut_lookup_le_miss_3_sva;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_2_nl = ~(lut_lookup_3_else_if_else_if_acc_itm_3_1
      | lut_lookup_else_if_lor_7_lpi_1_dfm_6);
  assign lut_lookup_else_mux_176_nl = MUX_s_1_2_2((lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_2_nl),
      lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2, lut_lookup_else_unequal_tmp_13);
  assign lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0 = MUX_s_1_2_2(lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2,
      (lut_lookup_else_mux_176_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_if_1_lut_lookup_if_1_and_13_nl = (lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[8])
      & (~ lut_lookup_if_1_lor_7_lpi_1_dfm_5);
  assign lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2((lut_lookup_if_1_lut_lookup_if_1_and_13_nl),
      lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2, lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6 = MUX_v_2_2_2((lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1[7:6]),
      (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13[7:6]), lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse = (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_mux_12_cse_mx0 = MUX_s_1_2_2(lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~(lut_lookup_le_miss_3_sva
      | lut_lookup_lo_miss_3_sva);
  assign lut_lookup_le_fraction_3_lpi_1_dfm_9 = lut_lookup_else_if_else_le_fra_3_sva_4
      & ({{34{lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2}},
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_6_land_3_lpi_1_dfm_7)) & ({{34{lut_lookup_3_else_if_else_if_acc_itm_3_1}},
      lut_lookup_3_else_if_else_if_acc_itm_3_1}) & (signext_35_1(~ lut_lookup_else_if_lor_7_lpi_1_dfm_6));
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = ({1'b1 ,
      (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_2_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2[8:0]),
      9'b111111111, (readslicef_248_1_247((lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl)))));
  assign lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_2_nl),
      9'b111111111, IsNaN_8U_23U_6_land_3_lpi_1_dfm_7));
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = ({1'b1
      , (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0];
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = readslicef_248_1_247((lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl));
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_2_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2[8:0]),
      9'b111111111, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1));
  assign lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_2_nl),
      9'b111111111, IsNaN_8U_23U_10_land_3_lpi_1_dfm_6));
  assign lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1 = (lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[7:0])
      & (signext_8_1(~ (lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[8]))) & (signext_8_1(~
      lut_lookup_if_1_lor_7_lpi_1_dfm_5));
  assign lut_lookup_lo_fraction_3_lpi_1_dfm_1 = lut_lookup_if_1_else_lo_fra_3_sva_4
      & ({{34{lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2}},
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_10_land_3_lpi_1_dfm_6)) & (signext_35_1(~ (lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[8])))
      & (signext_35_1(~ lut_lookup_if_1_lor_7_lpi_1_dfm_5));
  assign lut_lookup_3_else_2_and_svs = lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0
      & lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0;
  assign nl_lut_lookup_4_else_if_else_if_acc_nl = conv_u2u_3_4(lut_lookup_else_if_else_le_int_lpi_1_dfm_1[8:6])
      + 4'b1111;
  assign lut_lookup_4_else_if_else_if_acc_nl = nl_lut_lookup_4_else_if_else_if_acc_nl[3:0];
  assign lut_lookup_4_else_if_else_if_acc_itm_3_1 = readslicef_4_1_3((lut_lookup_4_else_if_else_if_acc_nl));
  assign lut_lookup_lo_miss_sva = lut_lookup_lo_uflow_lpi_1_dfm_4 | lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_sva = lut_lookup_le_uflow_lpi_1_dfm_6 | lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign lut_lookup_if_1_lut_lookup_if_1_and_14_nl = (lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[8])
      & (~ lut_lookup_if_1_lor_1_lpi_1_dfm_5);
  assign lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 = MUX_s_1_2_2((lut_lookup_if_1_lut_lookup_if_1_and_14_nl),
      lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2, lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse
      = lut_lookup_lo_miss_sva & lut_lookup_le_miss_sva;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_3_nl = ~(lut_lookup_4_else_if_else_if_acc_itm_3_1
      | lut_lookup_else_if_lor_1_lpi_1_dfm_6);
  assign lut_lookup_else_mux_178_nl = MUX_s_1_2_2((lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_3_nl),
      lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2, lut_lookup_else_unequal_tmp_13);
  assign lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0 = MUX_s_1_2_2(lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2,
      (lut_lookup_else_mux_178_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6 = MUX_v_2_2_2((lut_lookup_lo_index_0_7_0_lpi_1_dfm_1[7:6]),
      (lut_lookup_lo_index_0_7_0_lpi_1_dfm_13[7:6]), lut_lookup_unequal_tmp_13);
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse = (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_mux_17_cse_mx0 = MUX_s_1_2_2(lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~(lut_lookup_le_miss_sva
      | lut_lookup_lo_miss_sva);
  assign lut_lookup_le_fraction_lpi_1_dfm_9 = lut_lookup_else_if_else_le_fra_sva_4
      & ({{34{lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2}},
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_6_land_lpi_1_dfm_7)) & ({{34{lut_lookup_4_else_if_else_if_acc_itm_3_1}},
      lut_lookup_4_else_if_else_if_acc_itm_3_1}) & (signext_35_1(~ lut_lookup_else_if_lor_1_lpi_1_dfm_6));
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = ({1'b1 ,
      (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_3_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2[8:0]),
      9'b111111111, (readslicef_248_1_247((lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl)))));
  assign lut_lookup_else_if_else_le_int_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_3_nl),
      9'b111111111, IsNaN_8U_23U_6_land_lpi_1_dfm_7));
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = ({1'b1
      , (~ (FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2[255:9]))}) + 248'b1;
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0];
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = readslicef_248_1_247((lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl));
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_3_nl = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2[8:0]),
      9'b111111111, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1));
  assign lut_lookup_if_1_else_lo_int_lpi_1_dfm_1 = ~(MUX_v_9_2_2((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_3_nl),
      9'b111111111, IsNaN_8U_23U_10_land_lpi_1_dfm_6));
  assign lut_lookup_lo_index_0_7_0_lpi_1_dfm_1 = (lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[7:0])
      & (signext_8_1(~ (lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[8]))) & (signext_8_1(~
      lut_lookup_if_1_lor_1_lpi_1_dfm_5));
  assign lut_lookup_lo_fraction_lpi_1_dfm_1 = lut_lookup_if_1_else_lo_fra_sva_4 &
      ({{34{lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2}},
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2})
      & (signext_35_1(~ IsNaN_8U_23U_10_land_lpi_1_dfm_6)) & (signext_35_1(~ (lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[8])))
      & (signext_35_1(~ lut_lookup_if_1_lor_1_lpi_1_dfm_5));
  assign lut_lookup_4_else_2_and_svs = lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0 &
      lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0;
  assign lut_lookup_lut_lookup_nor_19_cse = ~(reg_lut_lookup_if_unequal_cse | cfg_lut_le_function_1_sva_10
      | lut_lookup_or_3_tmp);
  assign lut_lookup_and_5_cse = reg_lut_lookup_if_unequal_cse & (~ cfg_lut_le_function_1_sva_10)
      & (~ lut_lookup_or_3_tmp);
  assign lut_lookup_and_6_cse = (~ lut_lookup_unequal_tmp_13) & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_3_tmp);
  assign lut_lookup_and_7_cse = lut_lookup_unequal_tmp_13 & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_3_tmp);
  assign lut_lookup_or_3_tmp = (((lut_lookup_le_miss_1_sva & (~(lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse
      | lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs))) | (cfg_lut_hybrid_priority_1_sva_10
      & (lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse
      | lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs))) & (~(lut_lookup_1_else_2_and_svs
      | lut_lookup_1_and_svs_2))) | (cfg_lut_oflow_priority_1_sva_10 & lut_lookup_1_else_2_and_svs
      & (~ lut_lookup_1_and_svs_2)) | (cfg_lut_uflow_priority_1_sva_10 & lut_lookup_1_and_svs_2);
  assign lut_lookup_lut_lookup_nor_18_cse = ~(reg_lut_lookup_if_unequal_cse | cfg_lut_le_function_1_sva_10
      | lut_lookup_or_7_tmp);
  assign lut_lookup_and_13_cse = reg_lut_lookup_if_unequal_cse & (~ cfg_lut_le_function_1_sva_10)
      & (~ lut_lookup_or_7_tmp);
  assign lut_lookup_and_14_cse = (~ lut_lookup_else_unequal_tmp_13) & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_7_tmp);
  assign lut_lookup_and_15_cse = lut_lookup_else_unequal_tmp_13 & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_7_tmp);
  assign lut_lookup_or_7_tmp = (((lut_lookup_le_miss_2_sva & (~(lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse
      | lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs))) | (cfg_lut_hybrid_priority_1_sva_10
      & (lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse
      | lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs))) & (~(lut_lookup_2_else_2_and_svs
      | lut_lookup_2_and_svs_2))) | (cfg_lut_oflow_priority_1_sva_10 & lut_lookup_2_else_2_and_svs
      & (~ lut_lookup_2_and_svs_2)) | (cfg_lut_uflow_priority_1_sva_10 & lut_lookup_2_and_svs_2);
  assign lut_lookup_lut_lookup_nor_17_cse = ~(reg_lut_lookup_if_unequal_cse | cfg_lut_le_function_1_sva_10
      | lut_lookup_or_11_tmp);
  assign lut_lookup_and_21_cse = reg_lut_lookup_if_unequal_cse & (~ cfg_lut_le_function_1_sva_10)
      & (~ lut_lookup_or_11_tmp);
  assign lut_lookup_and_22_cse = (~ lut_lookup_else_unequal_tmp_13) & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_11_tmp);
  assign lut_lookup_and_23_cse = lut_lookup_else_unequal_tmp_13 & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_11_tmp);
  assign lut_lookup_or_11_tmp = (((lut_lookup_le_miss_3_sva & (~(lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse
      | lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs))) | (cfg_lut_hybrid_priority_1_sva_10
      & (lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse
      | lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs))) & (~(lut_lookup_3_else_2_and_svs
      | lut_lookup_3_and_svs_2))) | (cfg_lut_oflow_priority_1_sva_10 & lut_lookup_3_else_2_and_svs
      & (~ lut_lookup_3_and_svs_2)) | (cfg_lut_uflow_priority_1_sva_10 & lut_lookup_3_and_svs_2);
  assign lut_lookup_lut_lookup_nor_16_cse = ~(reg_lut_lookup_if_unequal_cse | cfg_lut_le_function_1_sva_10
      | lut_lookup_or_15_tmp);
  assign lut_lookup_and_29_cse = reg_lut_lookup_if_unequal_cse & (~ cfg_lut_le_function_1_sva_10)
      & (~ lut_lookup_or_15_tmp);
  assign lut_lookup_and_30_cse = (~ lut_lookup_else_unequal_tmp_13) & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_15_tmp);
  assign lut_lookup_and_31_cse = lut_lookup_else_unequal_tmp_13 & cfg_lut_le_function_1_sva_10
      & (~ lut_lookup_or_15_tmp);
  assign lut_lookup_or_15_tmp = (((lut_lookup_le_miss_sva & (~(lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse
      | lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs))) | (cfg_lut_hybrid_priority_1_sva_10
      & (lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse
      | lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs))) & (~(lut_lookup_4_else_2_and_svs
      | lut_lookup_4_and_svs_2))) | (cfg_lut_oflow_priority_1_sva_10 & lut_lookup_4_else_2_and_svs
      & (~ lut_lookup_4_and_svs_2)) | (cfg_lut_uflow_priority_1_sva_10 & lut_lookup_4_and_svs_2);
  assign main_stage_en_1 = chn_lut_in_rsci_bawt & or_cse;
  assign FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_19_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_1_sva, FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_1_sva,
      FpAdd_8U_23U_addend_larger_asn_19_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3,
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_30_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3,
      (FpAdd_8U_23U_is_a_greater_oelse_not_30_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_1_sva, FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_1_sva,
      FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1,
      FpAdd_8U_23U_2_a_int_mant_p1_1_sva, FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_a_int_mant_p1_1_sva,
      FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1, FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3,
      FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_is_a_greater_oelse_not_23_nl = ~ FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4;
  assign FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3,
      (FpAdd_8U_23U_2_is_a_greater_oelse_not_23_nl));
  assign FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_13_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_2_sva, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_2_sva,
      FpAdd_8U_23U_addend_larger_asn_13_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3,
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_32_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3,
      (FpAdd_8U_23U_is_a_greater_oelse_not_32_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_2_sva, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_2_sva,
      FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1,
      FpAdd_8U_23U_2_a_int_mant_p1_2_sva, FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_a_int_mant_p1_2_sva,
      FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1, FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3,
      FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_is_a_greater_oelse_not_25_nl = ~ FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4;
  assign FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3,
      (FpAdd_8U_23U_2_is_a_greater_oelse_not_25_nl));
  assign FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_7_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_3_sva, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_3_sva,
      FpAdd_8U_23U_addend_larger_asn_7_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3,
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_34_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3,
      (FpAdd_8U_23U_is_a_greater_oelse_not_34_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_3_sva, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_3_sva,
      FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1,
      FpAdd_8U_23U_2_a_int_mant_p1_3_sva, FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_a_int_mant_p1_3_sva,
      FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1, FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3,
      FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_is_a_greater_oelse_not_27_nl = ~ FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4;
  assign FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3,
      (FpAdd_8U_23U_2_is_a_greater_oelse_not_27_nl));
  assign FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_1_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_sva, FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_sva,
      FpAdd_8U_23U_addend_larger_asn_1_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_sva_3,
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_36_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_1_a_right_shift_qr_sva_3,
      (FpAdd_8U_23U_is_a_greater_oelse_not_36_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_sva, FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_sva,
      FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1,
      FpAdd_8U_23U_2_a_int_mant_p1_sva, FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_2_a_int_mant_p1_sva,
      FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1, FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_sva_3,
      FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_8U_23U_2_is_a_greater_oelse_not_29_nl = ~ FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4;
  assign FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, FpAdd_8U_23U_2_a_right_shift_qr_sva_3,
      (FpAdd_8U_23U_2_is_a_greater_oelse_not_29_nl));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_1_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_9);
  assign FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl),
      (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]);
  assign nl_lut_lookup_if_else_else_else_le_index_s_1_sva = conv_s2u_6_9({(reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[4:0]))}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_if_else_else_else_le_index_s_1_sva = nl_lut_lookup_if_else_else_else_le_index_s_1_sva[8:0];
  assign lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva = MUX_v_9_2_2((lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_1_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_itm, FpNormalize_8U_49U_2_oelse_not_9);
  assign FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_1_nl),
      (FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49:1]), FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49]);
  assign lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = MUX_v_9_2_2((lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_2_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_11);
  assign FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl),
      (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]);
  assign nl_lut_lookup_if_else_else_else_le_index_s_2_sva = conv_s2u_6_9({(reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[4:0]))}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_if_else_else_else_le_index_s_2_sva = nl_lut_lookup_if_else_else_else_le_index_s_2_sva[8:0];
  assign lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva = MUX_v_9_2_2((lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_3_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_itm, FpNormalize_8U_49U_2_oelse_not_11);
  assign FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_3_nl),
      (FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49:1]), FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49]);
  assign lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = MUX_v_9_2_2((lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_3_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_13);
  assign FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl),
      (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]);
  assign nl_lut_lookup_if_else_else_else_le_index_s_3_sva = conv_s2u_6_9({(reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[4:0]))}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_if_else_else_else_le_index_s_3_sva = nl_lut_lookup_if_else_else_else_le_index_s_3_sva[8:0];
  assign lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva = MUX_v_9_2_2((lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_5_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_itm, FpNormalize_8U_49U_2_oelse_not_13);
  assign FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_5_nl),
      (FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49:1]), FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49]);
  assign lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = MUX_v_9_2_2((lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_4_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_15);
  assign FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl),
      (FpAdd_8U_23U_1_int_mant_p1_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_sva_3[49]);
  assign nl_lut_lookup_if_else_else_else_le_index_s_sva = conv_s2u_6_9({(reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5])
      , (~ (reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[4:0]))}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_5);
  assign lut_lookup_if_else_else_else_le_index_s_sva = nl_lut_lookup_if_else_else_else_le_index_s_sva[8:0];
  assign lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva = MUX_v_9_2_2((lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl));
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_7_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_itm, FpNormalize_8U_49U_2_oelse_not_15);
  assign FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_7_nl),
      (FpAdd_8U_23U_2_int_mant_p1_sva_3[49:1]), FpAdd_8U_23U_2_int_mant_p1_sva_3[49]);
  assign lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136]!=151'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = MUX_v_9_2_2((lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127]),
      9'b111111111, (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl));
  assign nl_lut_lookup_1_if_if_else_else_if_acc_nl = conv_u2u_3_4(lut_lookup_if_if_else_else_le_index_s_1_sva[8:6])
      + 4'b1111;
  assign lut_lookup_1_if_if_else_else_if_acc_nl = nl_lut_lookup_1_if_if_else_else_if_acc_nl[3:0];
  assign lut_lookup_1_if_if_else_else_if_acc_itm_3 = readslicef_4_1_3((lut_lookup_1_if_if_else_else_if_acc_nl));
  assign nl_lut_lookup_if_if_else_else_le_index_s_1_sva = ({reg_lut_lookup_1_else_else_else_else_acc_reg
      , reg_lut_lookup_1_else_else_else_else_acc_1_reg , reg_lut_lookup_1_else_else_else_else_acc_2_reg
      , reg_lut_lookup_1_else_else_else_else_acc_3_reg}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_if_if_else_else_le_index_s_1_sva = nl_lut_lookup_if_if_else_else_le_index_s_1_sva[8:0];
  assign nl_lut_lookup_2_if_if_else_else_if_acc_nl = conv_u2u_3_4(lut_lookup_if_if_else_else_le_index_s_2_sva[8:6])
      + 4'b1111;
  assign lut_lookup_2_if_if_else_else_if_acc_nl = nl_lut_lookup_2_if_if_else_else_if_acc_nl[3:0];
  assign lut_lookup_2_if_if_else_else_if_acc_itm_3 = readslicef_4_1_3((lut_lookup_2_if_if_else_else_if_acc_nl));
  assign nl_lut_lookup_if_if_else_else_le_index_s_2_sva = ({reg_lut_lookup_2_else_else_else_else_acc_reg
      , reg_lut_lookup_2_else_else_else_else_acc_1_reg , reg_lut_lookup_2_else_else_else_else_acc_2_reg
      , reg_lut_lookup_2_else_else_else_else_acc_3_reg}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_if_if_else_else_le_index_s_2_sva = nl_lut_lookup_if_if_else_else_le_index_s_2_sva[8:0];
  assign nl_lut_lookup_3_if_if_else_else_if_acc_nl = conv_u2u_3_4(lut_lookup_if_if_else_else_le_index_s_3_sva[8:6])
      + 4'b1111;
  assign lut_lookup_3_if_if_else_else_if_acc_nl = nl_lut_lookup_3_if_if_else_else_if_acc_nl[3:0];
  assign lut_lookup_3_if_if_else_else_if_acc_itm_3 = readslicef_4_1_3((lut_lookup_3_if_if_else_else_if_acc_nl));
  assign nl_lut_lookup_if_if_else_else_le_index_s_3_sva = ({reg_lut_lookup_3_else_else_else_else_acc_reg
      , reg_lut_lookup_3_else_else_else_else_acc_1_reg , reg_lut_lookup_3_else_else_else_else_acc_2_reg
      , reg_lut_lookup_3_else_else_else_else_acc_3_reg}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_if_if_else_else_le_index_s_3_sva = nl_lut_lookup_if_if_else_else_le_index_s_3_sva[8:0];
  assign nl_lut_lookup_4_if_if_else_else_if_acc_nl = conv_u2u_3_4(lut_lookup_if_if_else_else_le_index_s_sva[8:6])
      + 4'b1111;
  assign lut_lookup_4_if_if_else_else_if_acc_nl = nl_lut_lookup_4_if_if_else_else_if_acc_nl[3:0];
  assign lut_lookup_4_if_if_else_else_if_acc_itm_3 = readslicef_4_1_3((lut_lookup_4_if_if_else_else_if_acc_nl));
  assign nl_lut_lookup_if_if_else_else_le_index_s_sva = ({reg_lut_lookup_4_else_else_else_else_acc_reg
      , reg_lut_lookup_4_else_else_else_else_acc_1_reg , reg_lut_lookup_4_else_else_else_else_acc_2_reg
      , reg_lut_lookup_4_else_else_else_else_acc_3_reg}) - conv_s2u_8_9(cfg_lut_le_index_offset_1_sva_7);
  assign lut_lookup_if_if_else_else_le_index_s_sva = nl_lut_lookup_if_if_else_else_le_index_s_sva[8:0];
  assign nl_lut_lookup_1_else_else_acc_1_nl = conv_s2u_32_33(cfg_lut_le_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[31:0]);
  assign lut_lookup_1_else_else_acc_1_nl = nl_lut_lookup_1_else_else_acc_1_nl[32:0];
  assign lut_lookup_1_else_else_acc_1_itm_32 = readslicef_33_1_32((lut_lookup_1_else_else_acc_1_nl));
  assign nl_lut_lookup_3_else_else_acc_1_nl = conv_s2u_32_33(cfg_lut_le_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[95:64]);
  assign lut_lookup_3_else_else_acc_1_nl = nl_lut_lookup_3_else_else_acc_1_nl[32:0];
  assign lut_lookup_3_else_else_acc_1_itm_32 = readslicef_33_1_32((lut_lookup_3_else_else_acc_1_nl));
  assign IsNaN_8U_23U_3_nor_4_tmp = ~((chn_lut_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_3_nor_6_tmp = ~((chn_lut_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000));
  assign nl_lut_lookup_2_else_else_acc_1_nl = conv_s2u_32_33(cfg_lut_le_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[63:32]);
  assign lut_lookup_2_else_else_acc_1_nl = nl_lut_lookup_2_else_else_acc_1_nl[32:0];
  assign lut_lookup_2_else_else_acc_1_itm_32 = readslicef_33_1_32((lut_lookup_2_else_else_acc_1_nl));
  assign IsNaN_8U_23U_3_nor_8_tmp = ~((chn_lut_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000));
  assign nl_lut_lookup_4_else_else_acc_1_nl = conv_s2u_32_33(cfg_lut_le_start_rsci_d)
      - conv_s2u_32_33(chn_lut_in_rsci_d_mxwt[127:96]);
  assign lut_lookup_4_else_else_acc_1_nl = nl_lut_lookup_4_else_else_acc_1_nl[32:0];
  assign lut_lookup_4_else_else_acc_1_itm_32 = readslicef_33_1_32((lut_lookup_4_else_else_acc_1_nl));
  assign IsNaN_8U_23U_3_nor_10_tmp = ~((chn_lut_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_4_nl = ({1'b1 , (cfg_lut_le_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[30:23])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_4_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_4_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_4_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_4_nl));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_6_nl = ({1'b1 , (cfg_lut_le_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[62:55])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_6_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_6_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_6_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_6_nl));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_8_nl = ({1'b1 , (cfg_lut_le_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[94:87])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_8_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_8_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_8_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_8_nl));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_10_nl = ({1'b1 , (cfg_lut_le_start_rsci_d[30:23])})
      + conv_u2u_8_9(~ (chn_lut_in_rsci_d_mxwt[126:119])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_10_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_10_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_10_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_10_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[22:0])})
      + conv_u2u_23_24(~ (cfg_lut_le_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[54:32])})
      + conv_u2u_23_24(~ (cfg_lut_le_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[86:64])})
      + conv_u2u_23_24(~ (cfg_lut_le_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[118:96])})
      + conv_u2u_23_24(~ (cfg_lut_le_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl));
  assign nl_lut_lookup_1_else_else_else_else_le_data_f_acc_2 = lut_lookup_1_else_else_else_else_le_data_f_lshift_1_itm
      + 32'b11111111111111111111111111111111;
  assign lut_lookup_1_else_else_else_else_le_data_f_acc_2 = nl_lut_lookup_1_else_else_else_else_le_data_f_acc_2[31:0];
  assign nl_lut_lookup_1_else_1_else_else_lo_data_f_acc_2 = lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_itm
      + 32'b11111111111111111111111111111111;
  assign lut_lookup_1_else_1_else_else_lo_data_f_acc_2 = nl_lut_lookup_1_else_1_else_else_lo_data_f_acc_2[31:0];
  assign nl_lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl = ({1'b1 , (~ reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm)
      , (~ reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm)}) + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)
      + 9'b1;
  assign lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl = nl_lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_9 = ((FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl)));
  assign nl_lut_lookup_1_FpNormalize_8U_49U_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)
      + 9'b1;
  assign lut_lookup_1_FpNormalize_8U_49U_2_acc_nl = nl_lut_lookup_1_FpNormalize_8U_49U_2_acc_nl[8:0];
  assign FpNormalize_8U_49U_2_oelse_not_9 = ((FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_1_FpNormalize_8U_49U_2_acc_nl)));
  assign nl_lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl = ({1'b1 , (~ reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm)
      , (~ reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm)}) + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)
      + 9'b1;
  assign lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl = nl_lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_11 = ((FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl)));
  assign nl_lut_lookup_2_FpNormalize_8U_49U_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)
      + 9'b1;
  assign lut_lookup_2_FpNormalize_8U_49U_2_acc_nl = nl_lut_lookup_2_FpNormalize_8U_49U_2_acc_nl[8:0];
  assign FpNormalize_8U_49U_2_oelse_not_11 = ((FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_2_FpNormalize_8U_49U_2_acc_nl)));
  assign nl_lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl = ({1'b1 , (~ reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm)
      , (~ reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm)}) + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16)
      + 9'b1;
  assign lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl = nl_lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_13 = ((FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl)));
  assign nl_lut_lookup_3_FpNormalize_8U_49U_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17)
      + 9'b1;
  assign lut_lookup_3_FpNormalize_8U_49U_2_acc_nl = nl_lut_lookup_3_FpNormalize_8U_49U_2_acc_nl[8:0];
  assign FpNormalize_8U_49U_2_oelse_not_13 = ((FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_3_FpNormalize_8U_49U_2_acc_nl)));
  assign nl_lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl = ({1'b1 , (~ reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm)
      , (~ reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm)}) + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18)
      + 9'b1;
  assign lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl = nl_lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_15 = ((FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl)));
  assign nl_lut_lookup_4_FpNormalize_8U_49U_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_qr_lpi_1_dfm_5)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19)
      + 9'b1;
  assign lut_lookup_4_FpNormalize_8U_49U_2_acc_nl = nl_lut_lookup_4_FpNormalize_8U_49U_2_acc_nl[8:0];
  assign FpNormalize_8U_49U_2_oelse_not_15 = ((FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((lut_lookup_4_FpNormalize_8U_49U_2_acc_nl)));
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm
      , (reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl = nl_lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0];
  assign lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = readslicef_8_1_7((lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl));
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm
      , (reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl = nl_lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0];
  assign lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = readslicef_8_1_7((lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl));
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm
      , (reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl = nl_lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0];
  assign lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = readslicef_8_1_7((lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl));
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm
      , (reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl = nl_lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0];
  assign lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = readslicef_8_1_7((lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl));
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm
      , (reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl = nl_lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0];
  assign lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl));
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm
      , (reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl = nl_lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0];
  assign lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl));
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm
      , (reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl = nl_lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0];
  assign lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl));
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl = ({1'b1 , reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm
      , (reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5:1])}) + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl = nl_lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0];
  assign lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl));
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp = ~((FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp!=8'b00000000));
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp = ~((FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7!=8'b00000000));
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp = ~((FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7!=8'b00000000));
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp = ~((FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0!=23'b00000000000000000000000)
      | (FpAdd_8U_23U_o_expo_lpi_1_dfm_7!=8'b00000000));
  assign or_tmp_6 = (~ chn_lut_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10);
  assign or_4_nl = nor_874_cse | (~ chn_lut_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10);
  assign mux_2_nl = MUX_s_1_2_2((~ main_stage_v_1), or_tmp_6, or_cse);
  assign mux_3_itm = MUX_s_1_2_2((mux_2_nl), (or_4_nl), or_26_cse);
  assign or_tmp_8 = (reg_cfg_precision_1_sva_st_12_cse_1[0]) | (~((reg_cfg_precision_1_sva_st_12_cse_1[1])
      & main_stage_v_1));
  assign mux_tmp_4 = MUX_s_1_2_2(or_1688_cse, or_tmp_6, or_cse);
  assign mux_tmp_10 = MUX_s_1_2_2(main_stage_v_2, main_stage_v_1, or_cse);
  assign nor_779_nl = ~((~ reg_chn_lut_out_rsci_ld_core_psct_cse) | chn_lut_out_rsci_bawt
      | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10));
  assign mux_18_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_1, or_cse);
  assign not_tmp_47 = MUX_s_1_2_2((mux_18_nl), (nor_779_nl), or_26_cse);
  assign mux_20_itm = MUX_s_1_2_2(or_1689_cse, or_tmp_8, or_cse);
  assign mux_25_itm = MUX_s_1_2_2(or_1689_cse, or_1688_cse, or_cse);
  assign or_tmp_44 = (reg_cfg_precision_1_sva_st_13_cse_1[0]) | (~((reg_cfg_precision_1_sva_st_13_cse_1[1])
      & main_stage_v_2));
  assign mux_26_itm = MUX_s_1_2_2(or_tmp_44, or_1688_cse, or_cse);
  assign mux_tmp_35 = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_cse);
  assign or_tmp_63 = (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10);
  assign and_tmp_5 = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & main_stage_v_3 & or_1857_cse;
  assign and_tmp_6 = main_stage_v_3 & or_1857_cse;
  assign or_tmp_101 = nor_13_cse | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10) |
      (~ main_stage_v_2);
  assign nor_tmp_12 = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 & lut_lookup_else_1_slc_32_mdf_1_sva_6
      & main_stage_v_2;
  assign nor_tmp_14 = lut_lookup_else_1_slc_32_mdf_1_sva_7 & FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign or_tmp_124 = (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10) | IsNaN_8U_23U_7_land_2_lpi_1_dfm_6
      | (~(IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 & main_stage_v_2));
  assign mux_70_nl = MUX_s_1_2_2(or_tmp_124, (~ main_stage_v_2), IsNaN_8U_23U_8_land_3_lpi_1_dfm_4);
  assign or_122_nl = (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10) | IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  assign mux_tmp_70 = MUX_s_1_2_2((mux_70_nl), or_tmp_124, or_122_nl);
  assign mux_72_nl = MUX_s_1_2_2(mux_tmp_70, (~ main_stage_v_2), IsNaN_8U_23U_8_land_1_lpi_1_dfm_6);
  assign or_121_nl = (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10) | IsNaN_8U_23U_7_land_1_lpi_1_dfm_6;
  assign mux_tmp_72 = MUX_s_1_2_2((mux_72_nl), mux_tmp_70, or_121_nl);
  assign or_tmp_129 = (cfg_precision_1_sva_st_70!=2'b10) | IsNaN_8U_23U_7_land_lpi_1_dfm_7
      | (~(IsNaN_8U_23U_8_land_lpi_1_dfm_5 & main_stage_v_3));
  assign mux_76_nl = MUX_s_1_2_2(or_tmp_129, (~ main_stage_v_3), IsNaN_8U_23U_8_land_3_lpi_1_dfm_5);
  assign or_127_nl = (cfg_precision_1_sva_st_70!=2'b10) | IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign mux_tmp_76 = MUX_s_1_2_2((mux_76_nl), or_tmp_129, or_127_nl);
  assign mux_78_nl = MUX_s_1_2_2(mux_tmp_76, (~ main_stage_v_3), IsNaN_8U_23U_8_land_2_lpi_1_dfm_7);
  assign or_126_nl = (cfg_precision_1_sva_st_70!=2'b10) | IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  assign mux_tmp_78 = MUX_s_1_2_2((mux_78_nl), mux_tmp_76, or_126_nl);
  assign nor_tmp_32 = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 & lut_lookup_else_1_slc_32_mdf_2_sva_6
      & main_stage_v_2;
  assign nor_tmp_34 = lut_lookup_else_1_slc_32_mdf_2_sva_7 & FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign nand_93_nl = ~(lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp & main_stage_v_2
      & (reg_cfg_precision_1_sva_st_13_cse_1==2'b10));
  assign or_191_nl = (~(lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49]))
      | lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp)) | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10);
  assign or_186_nl = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign mux_tmp_128 = MUX_s_1_2_2((or_191_nl), (nand_93_nl), or_186_nl);
  assign nand_tmp_4 = nor_874_cse | mux_tmp_128;
  assign and_tmp_14 = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & main_stage_v_3 & or_1857_cse;
  assign nor_tmp_44 = IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 & lut_lookup_else_1_slc_32_mdf_3_sva_6
      & main_stage_v_2;
  assign nor_tmp_46 = lut_lookup_else_1_slc_32_mdf_3_sva_7 & FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign and_tmp_19 = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & main_stage_v_3 & or_1857_cse;
  assign nor_tmp_55 = IsNaN_8U_23U_7_land_lpi_1_dfm_6 & lut_lookup_else_1_slc_32_mdf_sva_6
      & main_stage_v_2;
  assign nor_tmp_57 = lut_lookup_else_1_slc_32_mdf_sva_7 & FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign or_302_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 | IsNaN_8U_23U_8_land_lpi_1_dfm_5
      | IsNaN_8U_23U_7_land_lpi_1_dfm_7 | (cfg_precision_1_sva_st_70!=2'b10) | (~
      main_stage_v_3);
  assign mux_tmp_207 = MUX_s_1_2_2((or_302_nl), or_tmp_63, lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign or_tmp_314 = (cfg_precision_1_sva_st_71!=2'b10);
  assign not_tmp_209 = ~(lut_lookup_1_if_else_slc_32_svs_st_5 & main_stage_v_4 &
      or_tmp_314);
  assign mux_tmp_220 = MUX_s_1_2_2(main_stage_v_4, main_stage_v_3, or_cse);
  assign or_tmp_331 = FpAdd_8U_23U_2_mux_13_itm_3 | and_1141_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10);
  assign and_tmp_27 = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & main_stage_v_3 & or_1857_cse;
  assign not_tmp_222 = ~(lut_lookup_2_if_else_slc_32_svs_st_5 & main_stage_v_4 &
      or_tmp_314);
  assign or_tmp_363 = (cfg_precision_1_sva_st_70!=2'b10) | and_1140_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp
      | FpAdd_8U_23U_2_mux_29_itm_3 | (~ main_stage_v_3);
  assign not_tmp_235 = ~(lut_lookup_3_if_else_slc_32_svs_st_5 & main_stage_v_4 &
      or_tmp_314);
  assign or_tmp_378 = lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3 | not_tmp_235;
  assign or_tmp_380 = ~(cfg_lut_le_function_1_sva_st_42 & main_stage_v_4 & (cfg_precision_1_sva_st_71==2'b10));
  assign or_tmp_395 = FpAdd_8U_23U_2_mux_45_itm_3 | and_1139_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp
      | (cfg_precision_1_sva_st_70!=2'b10) | (~ main_stage_v_3);
  assign or_tmp_397 = lut_lookup_if_1_lor_7_lpi_1_dfm_4 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign not_tmp_248 = ~(lut_lookup_4_if_else_slc_32_svs_st_5 & main_stage_v_4 &
      or_tmp_314);
  assign or_tmp_427 = FpAdd_8U_23U_2_mux_61_itm_3 | and_1138_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp
      | (cfg_precision_1_sva_st_70!=2'b10) | (~ main_stage_v_3);
  assign or_tmp_428 = lut_lookup_if_1_lor_1_lpi_1_dfm_4 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_tmp_265 = MUX_s_1_2_2(main_stage_v_5, main_stage_v_4, or_cse);
  assign or_tmp_447 = ((lut_lookup_unequal_tmp_13 | (~ cfg_lut_le_function_1_sva_10))
      & lut_lookup_else_if_lor_5_lpi_1_dfm_6) | lut_lookup_else_if_lor_5_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse);
  assign mux_tmp_270 = MUX_s_1_2_2((~ main_stage_v_4), or_tmp_380, or_1853_cse);
  assign or_tmp_456 = (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse);
  assign mux_tmp_279 = IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 | lut_lookup_if_1_lor_5_lpi_1_dfm_4
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_tmp_281 = MUX_s_1_2_2((~ main_stage_v_4), or_312_cse, lut_lookup_else_unequal_tmp_18);
  assign or_tmp_478 = (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5);
  assign not_tmp_276 = ~((cfg_precision_1_sva_st_72[1]) & cfg_lut_le_function_1_sva_10
      & main_stage_v_5);
  assign mux_292_nl = MUX_s_1_2_2(or_tmp_380, (~ main_stage_v_4), cfg_lut_le_function_1_sva_st_42);
  assign mux_tmp_292 = MUX_s_1_2_2((mux_292_nl), or_tmp_380, lut_lookup_else_unequal_tmp_12);
  assign or_tmp_505 = (cfg_precision_1_sva_st_72[0]) | not_tmp_276;
  assign or_tmp_522 = (lut_lookup_unequal_tmp_13 & lut_lookup_if_1_lor_6_lpi_1_dfm_5)
      | lut_lookup_if_1_lor_6_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_107!=2'b10)
      | (~ main_stage_v_5);
  assign mux_tmp_301 = IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 | lut_lookup_if_1_lor_6_lpi_1_dfm_4
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign or_1851_cse = lut_lookup_else_unequal_tmp_13 | (~ cfg_lut_le_function_1_sva_10);
  assign or_tmp_547 = (or_1851_cse & lut_lookup_else_if_lor_7_lpi_1_dfm_6) | lut_lookup_else_if_lor_7_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse);
  assign and_850_cse = lut_lookup_unequal_tmp_13 & lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  assign or_tmp_573 = IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 | lut_lookup_if_1_lor_7_lpi_1_dfm_4
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign or_tmp_598 = (or_1851_cse & lut_lookup_else_if_lor_1_lpi_1_dfm_6) | lut_lookup_else_if_lor_1_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse);
  assign and_848_cse = lut_lookup_unequal_tmp_13 & lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign or_tmp_623 = IsNaN_8U_23U_10_land_lpi_1_dfm_5 | lut_lookup_if_1_lor_1_lpi_1_dfm_4
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign not_tmp_334 = ~(cfg_lut_le_function_1_sva_10 | (~ main_stage_v_5));
  assign nor_tmp_112 = lut_lookup_else_unequal_tmp_18 & main_stage_v_4;
  assign mux_tmp_475 = MUX_s_1_2_2(or_1689_cse, (~ or_1689_cse), nor_42_cse);
  assign not_tmp_394 = ~((reg_cfg_precision_1_sva_st_12_cse_1[1]) | (~ mux_tmp_475));
  assign not_tmp_412 = ~((reg_cfg_precision_1_sva_st_12_cse_1[1]) | or_1689_cse);
  assign not_tmp_418 = ~((reg_cfg_precision_1_sva_st_12_cse_1[1]) | (~ or_1689_cse));
  assign not_tmp_422 = ~((reg_cfg_precision_1_sva_st_12_cse_1[1]) | (~ main_stage_v_1));
  assign nand_95_cse = ~(main_stage_v_1 & (reg_cfg_precision_1_sva_st_12_cse_1==2'b10));
  assign mux_581_nl = MUX_s_1_2_2(or_1688_cse, nand_95_cse, reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse);
  assign mux_582_itm = MUX_s_1_2_2((mux_581_nl), or_tmp_6, or_cse);
  assign mux_594_nl = MUX_s_1_2_2(or_1688_cse, nand_95_cse, reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse);
  assign mux_595_itm = MUX_s_1_2_2((mux_594_nl), or_tmp_6, or_cse);
  assign mux_tmp_595 = MUX_s_1_2_2(or_1689_cse, (~ or_1689_cse), nor_13_cse);
  assign or_1860_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4
      | (~ main_stage_v_1) | mux_tmp_595;
  assign mux_tmp_596 = MUX_s_1_2_2(mux_tmp_595, (or_1860_nl), nor_648_cse);
  assign or_tmp_843 = (cfg_precision_rsci_d!=2'b10) | (~(chn_lut_in_rsci_bawt & or_cse));
  assign mux_615_nl = MUX_s_1_2_2(or_tmp_843, (~ or_cse), FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49]);
  assign mux_616_nl = MUX_s_1_2_2((mux_615_nl), or_tmp_843, lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1);
  assign mux_617_nl = MUX_s_1_2_2((~ or_tmp_843), (~ (mux_616_nl)), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign or_841_nl = (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign mux_tmp_617 = MUX_s_1_2_2((mux_617_nl), (~ or_tmp_843), or_841_nl);
  assign nor_647_nl = ~(lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 | (~((FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49])
      & or_cse)));
  assign or_832_nl = IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  assign mux_tmp_618 = MUX_s_1_2_2((nor_647_nl), mux_tmp_617, or_832_nl);
  assign or_856_nl = IsNaN_8U_23U_7_land_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  assign mux_639_nl = MUX_s_1_2_2((~ main_stage_v_2), or_1689_cse, or_856_nl);
  assign mux_tmp_643 = MUX_s_1_2_2(or_1689_cse, (mux_639_nl), nor_196_cse);
  assign and_tmp_59 = reg_cfg_lut_le_function_1_sva_st_20_cse & IsNaN_8U_23U_1_land_1_lpi_1_dfm_7
      & main_stage_v_2 & or_66_cse;
  assign and_tmp_61 = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 & or_66_cse & main_stage_v_2;
  assign nor_641_nl = ~((reg_cfg_precision_1_sva_st_13_cse_1[1]) | (~ main_stage_v_2));
  assign mux_tmp_655 = MUX_s_1_2_2((nor_641_nl), main_stage_v_2, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign and_tmp_69 = IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 & main_stage_v_2 & or_66_cse;
  assign nor_622_nl = ~((cfg_precision_1_sva_st_70[1]) | (~ main_stage_v_3));
  assign mux_tmp_704 = MUX_s_1_2_2((nor_622_nl), main_stage_v_3, cfg_precision_1_sva_st_70[0]);
  assign and_tmp_83 = main_stage_v_4 & or_tmp_314;
  assign or_tmp_976 = (cfg_precision_1_sva_st_70!=2'b10) | cfg_lut_le_function_1_sva_st_41
      | (~ main_stage_v_3);
  assign or_tmp_980 = (cfg_precision_1_sva_8!=2'b10) | cfg_lut_le_function_1_sva_st_42
      | (~ main_stage_v_4);
  assign or_tmp_993 = nor_610_cse | cfg_lut_le_function_1_sva_st_42 | (~ main_stage_v_4);
  assign and_tmp_92 = lut_lookup_else_else_else_asn_mdf_1_sva_3 & cfg_lut_le_function_1_sva_st_41
      & FpAdd_8U_23U_1_mux_13_itm_4 & lut_lookup_else_else_slc_32_mdf_1_sva_7 & FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6
      & main_stage_v_3 & or_1857_cse;
  assign nor_tmp_238 = cfg_lut_le_function_1_sva_st_42 & IsNaN_8U_23U_6_land_1_lpi_1_dfm_6
      & lut_lookup_else_else_slc_32_mdf_1_sva_8 & main_stage_v_4;
  assign mux_793_cse = MUX_s_1_2_2(main_stage_v_3, and_tmp_6, nor_792_cse);
  assign and_tmp_97 = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 & lut_lookup_else_1_slc_32_mdf_1_sva_7
      & main_stage_v_3 & or_1857_cse;
  assign or_tmp_1043 = FpMantRNE_49U_24U_2_else_carry_1_sva_2 | FpAdd_8U_23U_2_mux_13_itm_3
      | (~ and_tmp_97);
  assign and_tmp_98 = lut_lookup_else_1_slc_32_mdf_1_sva_8 & IsNaN_8U_23U_10_land_1_lpi_1_dfm_5
      & main_stage_v_4 & or_tmp_314;
  assign and_tmp_103 = lut_lookup_else_else_else_asn_mdf_2_sva_3 & cfg_lut_le_function_1_sva_st_41
      & FpAdd_8U_23U_1_mux_29_itm_4 & FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & lut_lookup_else_else_slc_32_mdf_2_sva_7
      & main_stage_v_3 & or_1857_cse;
  assign nor_tmp_260 = cfg_lut_le_function_1_sva_st_42 & IsNaN_8U_23U_6_land_2_lpi_1_dfm_6
      & lut_lookup_else_else_slc_32_mdf_2_sva_8 & main_stage_v_4;
  assign nand_tmp_22 = ~(FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 & (~(nor_792_cse | FpMantRNE_49U_24U_2_else_carry_2_sva_2
      | FpAdd_8U_23U_2_mux_29_itm_3 | (~(lut_lookup_else_1_slc_32_mdf_2_sva_7 & main_stage_v_3)))));
  assign and_tmp_108 = lut_lookup_else_1_slc_32_mdf_2_sva_8 & IsNaN_8U_23U_10_land_2_lpi_1_dfm_5
      & main_stage_v_4 & or_tmp_314;
  assign and_tmp_113 = lut_lookup_else_else_else_asn_mdf_3_sva_3 & cfg_lut_le_function_1_sva_st_41
      & FpAdd_8U_23U_1_mux_45_itm_4 & lut_lookup_else_else_slc_32_mdf_3_sva_7 & FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6
      & main_stage_v_3 & or_1857_cse;
  assign nor_tmp_281 = cfg_lut_le_function_1_sva_st_42 & IsNaN_8U_23U_6_land_3_lpi_1_dfm_6
      & lut_lookup_else_else_slc_32_mdf_3_sva_8 & main_stage_v_4;
  assign or_tmp_1181 = FpAdd_8U_23U_2_mux_45_itm_3 | (~ FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5)
      | FpMantRNE_49U_24U_2_else_carry_3_sva_2 | (~(lut_lookup_else_1_slc_32_mdf_3_sva_7
      & and_tmp_6));
  assign and_tmp_119 = lut_lookup_else_1_slc_32_mdf_3_sva_8 & IsNaN_8U_23U_10_land_3_lpi_1_dfm_5
      & main_stage_v_4 & or_tmp_314;
  assign and_tmp_124 = lut_lookup_else_else_else_asn_mdf_sva_3 & cfg_lut_le_function_1_sva_st_41
      & FpAdd_8U_23U_1_mux_61_itm_4 & FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & lut_lookup_else_else_slc_32_mdf_sva_7
      & main_stage_v_3 & or_1857_cse;
  assign and_tmp_130 = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 & lut_lookup_else_1_slc_32_mdf_sva_7
      & and_tmp_6;
  assign or_tmp_1250 = FpMantRNE_49U_24U_2_else_carry_sva_2 | FpAdd_8U_23U_2_mux_61_itm_3
      | (~ and_tmp_130);
  assign and_tmp_131 = lut_lookup_else_1_slc_32_mdf_sva_8 & IsNaN_8U_23U_10_land_lpi_1_dfm_5
      & main_stage_v_4 & or_tmp_314;
  assign mux_tmp_978 = MUX_s_1_2_2(and_852_cse, and_826_cse, or_cse);
  assign or_tmp_1360 = and_794_cse | (~ chn_lut_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10);
  assign not_tmp_800 = ~(lut_lookup_1_if_else_slc_32_svs_6 & IsNaN_8U_23U_1_land_1_lpi_1_dfm_7
      & main_stage_v_2 & or_66_cse);
  assign or_tmp_1450 = (~ reg_chn_lut_out_rsci_ld_core_psct_cse) | chn_lut_out_rsci_bawt
      | reg_cfg_lut_le_function_1_sva_st_20_cse | not_tmp_800;
  assign mux_tmp_1101 = MUX_s_1_2_2(not_tmp_422, main_stage_v_1, or_26_cse);
  assign mux_tmp_1104 = main_stage_v_1 & or_26_cse;
  assign or_1495_cse = (cfg_precision_rsci_d!=2'b10);
  assign and_tmp_178 = chn_lut_in_rsci_bawt & or_1495_cse;
  assign and_dcpl_54 = (~ chn_lut_out_rsci_bawt) & reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign and_dcpl_59 = or_cse & main_stage_v_5 & (~ lut_lookup_1_and_svs_2);
  assign and_dcpl_63 = or_cse & main_stage_v_5 & (~ lut_lookup_2_and_svs_2);
  assign and_dcpl_67 = or_cse & main_stage_v_5 & (~ lut_lookup_3_and_svs_2);
  assign and_dcpl_71 = or_cse & main_stage_v_5 & (~ lut_lookup_4_and_svs_2);
  assign and_dcpl_72 = or_cse & main_stage_v_5;
  assign and_dcpl_74 = (~ main_stage_v_5) & chn_lut_out_rsci_bawt & reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign or_tmp_1490 = (~ reg_chn_lut_out_rsci_ld_core_psct_cse) | chn_lut_out_rsci_bawt
      | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10);
  assign and_dcpl_98 = (reg_cfg_precision_1_sva_st_13_cse_1==2'b10);
  assign and_dcpl_148 = or_cse & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign or_dcpl_51 = (~ or_66_cse) | reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign and_dcpl_161 = or_66_cse & or_cse;
  assign and_dcpl_162 = or_cse & (~ reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign or_dcpl_57 = and_dcpl_98 | reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign or_1583_nl = lut_lookup_if_if_lor_5_lpi_1_dfm_4 | (~((~ lut_lookup_1_if_if_else_acc_itm_9_1)
      | IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 | (cfg_precision_1_sva_st_71!=2'b10)));
  assign mux_1129_nl = MUX_s_1_2_2(lut_lookup_if_else_lut_lookup_if_else_or_cse,
      (or_1583_nl), nor_610_cse);
  assign mux_tmp_1130 = MUX_s_1_2_2((mux_1129_nl), lut_lookup_else_mux_itm_2, cfg_lut_le_function_1_sva_st_42);
  assign or_tmp_1513 = lut_lookup_lo_uflow_1_lpi_1_dfm_3 | mux_tmp_1130;
  assign mux_tmp_1136 = MUX_s_1_2_2((~ mux_tmp_1130), mux_tmp_1130, lut_lookup_lo_uflow_1_lpi_1_dfm_3);
  assign or_1594_nl = lut_lookup_if_if_lor_6_lpi_1_dfm_4 | (~((~ lut_lookup_2_if_if_else_acc_itm_9_1)
      | IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 | (cfg_precision_1_sva_st_71!=2'b10)));
  assign mux_1142_nl = MUX_s_1_2_2(lut_lookup_if_else_lut_lookup_if_else_or_1_cse,
      (or_1594_nl), nor_610_cse);
  assign mux_tmp_1143 = MUX_s_1_2_2((mux_1142_nl), lut_lookup_else_mux_43_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign or_tmp_1523 = lut_lookup_lo_uflow_2_lpi_1_dfm_3 | mux_tmp_1143;
  assign mux_tmp_1149 = MUX_s_1_2_2((~ mux_tmp_1143), mux_tmp_1143, lut_lookup_lo_uflow_2_lpi_1_dfm_3);
  assign or_1606_nl = lut_lookup_if_if_lor_7_lpi_1_dfm_4 | (~((~ lut_lookup_3_if_if_else_acc_itm_9_1)
      | IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 | (cfg_precision_1_sva_st_71!=2'b10)));
  assign mux_1155_nl = MUX_s_1_2_2(lut_lookup_if_else_lut_lookup_if_else_or_2_cse,
      (or_1606_nl), nor_610_cse);
  assign mux_tmp_1156 = MUX_s_1_2_2((mux_1155_nl), lut_lookup_else_mux_86_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign or_tmp_1534 = lut_lookup_lo_uflow_3_lpi_1_dfm_3 | mux_tmp_1156;
  assign mux_tmp_1162 = MUX_s_1_2_2((~ mux_tmp_1156), mux_tmp_1156, lut_lookup_lo_uflow_3_lpi_1_dfm_3);
  assign or_1618_nl = lut_lookup_if_if_lor_1_lpi_1_dfm_4 | (~((~ lut_lookup_4_if_if_else_acc_itm_9_1)
      | IsNaN_8U_23U_6_land_lpi_1_dfm_6 | (cfg_precision_1_sva_st_71!=2'b10)));
  assign mux_1168_nl = MUX_s_1_2_2(lut_lookup_if_else_lut_lookup_if_else_or_3_cse,
      (or_1618_nl), nor_610_cse);
  assign mux_tmp_1169 = MUX_s_1_2_2((mux_1168_nl), lut_lookup_else_mux_129_itm_2,
      cfg_lut_le_function_1_sva_st_42);
  assign or_tmp_1545 = lut_lookup_lo_uflow_lpi_1_dfm_3 | mux_tmp_1169;
  assign mux_tmp_1175 = MUX_s_1_2_2((~ mux_tmp_1169), mux_tmp_1169, lut_lookup_lo_uflow_lpi_1_dfm_3);
  assign and_dcpl_258 = or_cse & cfg_lut_le_function_1_sva_st_42;
  assign and_dcpl_259 = or_cse & (~ cfg_lut_le_function_1_sva_st_42);
  assign and_dcpl_280 = or_cse & (~ FpAdd_8U_23U_1_is_a_greater_acc_4_itm_8_1) &
      ((~ lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1);
  assign and_dcpl_284 = or_cse & ((~ lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_itm_23_1) & (~ FpAdd_8U_23U_2_is_a_greater_acc_itm_8_1);
  assign and_dcpl_288 = or_cse & ((~ lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1) & (~ FpAdd_8U_23U_1_is_a_greater_acc_6_itm_8_1);
  assign and_dcpl_292 = or_cse & ((~ lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_itm_23_1) & (~ FpAdd_8U_23U_2_is_a_greater_acc_1_itm_8_1);
  assign and_dcpl_296 = or_cse & ((~ lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1) & (~ FpAdd_8U_23U_1_is_a_greater_acc_8_itm_8_1);
  assign and_dcpl_300 = or_cse & ((~ lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_itm_23_1) & (~ FpAdd_8U_23U_2_is_a_greater_acc_2_itm_8_1);
  assign and_dcpl_304 = or_cse & (~ FpAdd_8U_23U_1_is_a_greater_acc_10_itm_8_1) &
      ((~ lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1);
  assign and_dcpl_308 = or_cse & ((~ lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_itm_23_1) & (~ FpAdd_8U_23U_2_is_a_greater_acc_3_itm_8_1);
  assign and_dcpl_309 = (cfg_precision_rsci_d==2'b10);
  assign and_dcpl_314 = or_1495_cse & or_cse;
  assign and_dcpl_315 = or_cse & cfg_lut_le_function_rsci_d;
  assign and_dcpl_316 = or_cse & (~ cfg_lut_le_function_rsci_d);
  assign and_dcpl_351 = or_cse & (~ (reg_cfg_precision_1_sva_st_12_cse_1[0]));
  assign and_dcpl_364 = and_956_cse & main_stage_v_1;
  assign and_dcpl_403 = or_1857_cse & cfg_lut_le_function_1_sva_st_41 & or_cse;
  assign and_dcpl_405 = and_896_cse & (~ cfg_lut_le_function_1_sva_st_41) & or_cse;
  assign or_tmp_1628 = or_cse & chn_lut_in_rsci_bawt & (fsm_output[1]);
  assign chn_lut_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign main_stage_v_1_mx0c1 = main_stage_v_1 & (~ chn_lut_in_rsci_bawt) & or_cse;
  assign main_stage_v_2_mx0c1 = main_stage_v_2 & (~ main_stage_v_1) & or_cse;
  assign main_stage_v_3_mx0c1 = main_stage_v_3 & (~ main_stage_v_2) & or_cse;
  assign main_stage_v_4_mx0c1 = (~ main_stage_v_3) & main_stage_v_4 & or_cse;
  assign main_stage_v_5_mx0c1 = main_stage_v_5 & (~ main_stage_v_4) & or_cse;
  assign nor_444_nl = ~(cfg_lut_uflow_priority_1_sva_9 | (~(lut_lookup_lo_uflow_1_lpi_1_dfm_3
      & mux_tmp_1130)));
  assign mux_1140_nl = MUX_s_1_2_2(or_tmp_1513, (~ mux_tmp_1136), cfg_lut_uflow_priority_1_sva_9);
  assign mux_1141_nl = MUX_s_1_2_2((mux_1140_nl), (nor_444_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1 = (mux_1141_nl) & or_cse;
  assign nor_442_nl = ~(cfg_lut_uflow_priority_1_sva_9 | (~(lut_lookup_lo_uflow_2_lpi_1_dfm_3
      & mux_tmp_1143)));
  assign mux_1153_nl = MUX_s_1_2_2(or_tmp_1523, (~ mux_tmp_1149), cfg_lut_uflow_priority_1_sva_9);
  assign mux_1154_nl = MUX_s_1_2_2((mux_1153_nl), (nor_442_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1 = (mux_1154_nl) & or_cse;
  assign nor_440_nl = ~(cfg_lut_uflow_priority_1_sva_9 | (~(lut_lookup_lo_uflow_3_lpi_1_dfm_3
      & mux_tmp_1156)));
  assign mux_1166_nl = MUX_s_1_2_2(or_tmp_1534, (~ mux_tmp_1162), cfg_lut_uflow_priority_1_sva_9);
  assign mux_1167_nl = MUX_s_1_2_2((mux_1166_nl), (nor_440_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1 = (mux_1167_nl) & or_cse;
  assign nor_438_nl = ~(cfg_lut_uflow_priority_1_sva_9 | (~(lut_lookup_lo_uflow_lpi_1_dfm_3
      & mux_tmp_1169)));
  assign mux_1179_nl = MUX_s_1_2_2(or_tmp_1545, (~ mux_tmp_1175), cfg_lut_uflow_priority_1_sva_9);
  assign mux_1180_nl = MUX_s_1_2_2((mux_1179_nl), (nor_438_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1 = (mux_1180_nl) & or_cse;
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[22:0])})
      + conv_u2u_23_24(~ (cfg_lut_lo_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl[23:0];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[54:32])})
      + conv_u2u_23_24(~ (cfg_lut_lo_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl[23:0];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[86:64])})
      + conv_u2u_23_24(~ (cfg_lut_lo_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl[23:0];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , (chn_lut_in_rsci_d_mxwt[118:96])})
      + conv_u2u_23_24(~ (cfg_lut_lo_start_rsci_d[22:0])) + 24'b1;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl[23:0];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl));
  assign nl_lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = nl_lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = nl_lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = nl_lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = nl_lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = nl_lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = nl_lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = nl_lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = nl_lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0];
  assign and_553_m1c = or_cse & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_6) & reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_555_m1c = or_cse & (~(IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 | reg_cfg_lut_le_function_1_sva_st_19_cse));
  assign and_590_m1c = reg_cfg_lut_le_function_1_sva_st_19_cse & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_6)
      & or_cse;
  assign and_592_m1c = (~(reg_cfg_lut_le_function_1_sva_st_19_cse | reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse))
      & or_cse;
  assign chn_lut_in_rsci_oswt_unreg = or_tmp_1628;
  assign chn_lut_out_rsci_oswt_unreg = chn_lut_out_rsci_bawt & reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign and_dcpl_540 = core_wen & main_stage_v_1;
  assign or_tmp_1663 = nor_193_cse | (~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_1_if_else_else_acc_itm_10 | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7);
  assign and_dcpl_576 = main_stage_v_2 & core_wen;
  assign or_tmp_1671 = (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7) | reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign or_tmp_1674 = nor_193_cse | (~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_2_if_else_else_acc_itm_10 | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7);
  assign or_tmp_1678 = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_2_if_else_else_acc_itm_10;
  assign or_tmp_1684 = nor_193_cse | (~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_3_if_else_else_acc_itm_10 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7);
  assign or_1972_nl = IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 | nor_38_cse_1;
  assign or_1973_nl = IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 | nor_38_cse_1;
  assign mux_1234_nl = MUX_s_1_2_2((or_1973_nl), (or_1972_nl), reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign or_tmp_1692 = lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp | (~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      | (mux_1234_nl)));
  assign or_tmp_1697 = nor_193_cse | (~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_4_if_else_else_acc_itm_10 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7);
  assign or_1991_nl = IsNaN_8U_23U_4_land_lpi_1_dfm_4 | nor_50_cse_1;
  assign or_1992_nl = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse | nor_50_cse_1;
  assign mux_1241_nl = MUX_s_1_2_2((or_1992_nl), (or_1991_nl), reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign or_tmp_1705 = lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp | (~(IsNaN_8U_23U_1_land_lpi_1_dfm_7
      | (mux_1241_nl)));
  assign or_tmp_1707 = (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7) | reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign and_dcpl_648 = core_wen & main_stage_v_3;
  assign or_tmp_1716 = (~ FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_1_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_1_sva_7);
  assign or_tmp_1720 = nor_792_cse | (~ FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_2_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_2_sva_7);
  assign nor_823_nl = ~((~((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2[8])
      | lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1)) | lut_lookup_if_1_lor_5_lpi_1_dfm_5
      | IsNaN_8U_23U_10_land_1_lpi_1_dfm_6);
  assign mux_tmp_1247 = MUX_s_1_2_2((nor_823_nl), lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2,
      lut_lookup_unequal_tmp_13);
  assign nor_820_nl = ~(lut_lookup_if_1_lor_6_lpi_1_dfm_5 | (~((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2[8])
      | lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1)) | IsNaN_8U_23U_10_land_2_lpi_1_dfm_6);
  assign mux_tmp_1250 = MUX_s_1_2_2((nor_820_nl), lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2,
      lut_lookup_unequal_tmp_13);
  assign nor_817_nl = ~((~((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2[8])
      | lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1)) | lut_lookup_if_1_lor_7_lpi_1_dfm_5
      | IsNaN_8U_23U_10_land_3_lpi_1_dfm_6);
  assign mux_tmp_1253 = MUX_s_1_2_2((nor_817_nl), lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2,
      lut_lookup_unequal_tmp_13);
  assign nor_813_cse = ~((FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2[8]) | lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1);
  assign or_2056_nl = lut_lookup_unequal_tmp_13 | (~ IsNaN_8U_23U_10_land_lpi_1_dfm_6);
  assign or_2055_nl = nor_813_cse | lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign mux_1261_nl = MUX_s_1_2_2((or_2056_nl), lut_lookup_unequal_tmp_13, or_2055_nl);
  assign nor_814_nl = ~(nor_813_cse | lut_lookup_if_1_lor_1_lpi_1_dfm_5 | lut_lookup_unequal_tmp_13
      | IsNaN_8U_23U_10_land_lpi_1_dfm_6);
  assign mux_tmp_1257 = MUX_s_1_2_2((nor_814_nl), (mux_1261_nl), lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2);
  assign and_tmp_201 = lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 & mux_tmp_1257;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp = (fsm_output[1]) & FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp = (fsm_output[1]) & FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1 = (fsm_output[1]) & FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp_1 = (fsm_output[1]) & FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp_2 = (fsm_output[1]) & FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2 = (fsm_output[1]) & FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3 = (fsm_output[1]) & FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp_3 = (fsm_output[1]) & FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_in_rsci_iswt0 <= 1'b0;
      chn_lut_out_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_lut_in_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_lut_out_rsci_iswt0 <= and_dcpl_72;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_lut_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_lut_in_rsci_ld_core_psct <= chn_lut_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_d_11_0 <= 12'b0;
      chn_lut_out_rsci_d_34_12 <= 23'b0;
      chn_lut_out_rsci_d_46_35 <= 12'b0;
      chn_lut_out_rsci_d_69_47 <= 23'b0;
      chn_lut_out_rsci_d_81_70 <= 12'b0;
      chn_lut_out_rsci_d_104_82 <= 23'b0;
      chn_lut_out_rsci_d_116_105 <= 12'b0;
      chn_lut_out_rsci_d_139_117 <= 23'b0;
      chn_lut_out_rsci_d_267_140 <= 128'b0;
      chn_lut_out_rsci_d_268 <= 1'b0;
      chn_lut_out_rsci_d_269 <= 1'b0;
      chn_lut_out_rsci_d_270 <= 1'b0;
      chn_lut_out_rsci_d_271 <= 1'b0;
      chn_lut_out_rsci_d_285_280 <= 6'b0;
      chn_lut_out_rsci_d_294_289 <= 6'b0;
      chn_lut_out_rsci_d_303_298 <= 6'b0;
      chn_lut_out_rsci_d_312_307 <= 6'b0;
      chn_lut_out_rsci_d_316 <= 1'b0;
      chn_lut_out_rsci_d_317 <= 1'b0;
      chn_lut_out_rsci_d_318 <= 1'b0;
      chn_lut_out_rsci_d_319 <= 1'b0;
      chn_lut_out_rsci_d_320 <= 1'b0;
      chn_lut_out_rsci_d_321 <= 1'b0;
      chn_lut_out_rsci_d_322 <= 1'b0;
      chn_lut_out_rsci_d_323 <= 1'b0;
    end
    else if ( chn_lut_out_and_cse ) begin
      chn_lut_out_rsci_d_11_0 <= MUX_v_12_2_2(12'b000000000000, (lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_7_nl),
          (lut_lookup_not_39_nl));
      chn_lut_out_rsci_d_34_12 <= MUX1HOT_v_23_6_2(lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1,
          (lut_lookup_le_fraction_1_lpi_1_dfm_22[34:12]), (lut_lookup_le_fraction_1_lpi_1_dfm_9[34:12]),
          (lut_lookup_le_fraction_1_lpi_1_dfm_21[34:12]), (lut_lookup_lo_fraction_1_lpi_1_dfm_1[34:12]),
          (lut_lookup_lo_fraction_1_lpi_1_dfm_9[34:12]), {lut_lookup_lut_lookup_nor_19_cse
          , lut_lookup_and_5_cse , lut_lookup_and_6_cse , lut_lookup_and_7_cse ,
          lut_lookup_and_138_cse , lut_lookup_and_139_cse});
      chn_lut_out_rsci_d_46_35 <= MUX_v_12_2_2(12'b000000000000, (lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_6_nl),
          (lut_lookup_not_38_nl));
      chn_lut_out_rsci_d_69_47 <= MUX1HOT_v_23_6_2(lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1,
          (lut_lookup_le_fraction_2_lpi_1_dfm_22[34:12]), (lut_lookup_le_fraction_2_lpi_1_dfm_9[34:12]),
          (lut_lookup_le_fraction_2_lpi_1_dfm_21[34:12]), (lut_lookup_lo_fraction_2_lpi_1_dfm_1[34:12]),
          (lut_lookup_lo_fraction_2_lpi_1_dfm_9[34:12]), {lut_lookup_lut_lookup_nor_18_cse
          , lut_lookup_and_13_cse , lut_lookup_and_14_cse , lut_lookup_and_15_cse
          , lut_lookup_and_136_cse , lut_lookup_and_137_cse});
      chn_lut_out_rsci_d_81_70 <= MUX_v_12_2_2(12'b000000000000, (lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_5_nl),
          (lut_lookup_not_37_nl));
      chn_lut_out_rsci_d_104_82 <= MUX1HOT_v_23_6_2(lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1,
          (lut_lookup_le_fraction_3_lpi_1_dfm_22[34:12]), (lut_lookup_le_fraction_3_lpi_1_dfm_9[34:12]),
          (lut_lookup_le_fraction_3_lpi_1_dfm_21[34:12]), (lut_lookup_lo_fraction_3_lpi_1_dfm_1[34:12]),
          (lut_lookup_lo_fraction_3_lpi_1_dfm_9[34:12]), {lut_lookup_lut_lookup_nor_17_cse
          , lut_lookup_and_21_cse , lut_lookup_and_22_cse , lut_lookup_and_23_cse
          , lut_lookup_and_134_cse , lut_lookup_and_135_cse});
      chn_lut_out_rsci_d_116_105 <= MUX_v_12_2_2(12'b000000000000, (lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_4_nl),
          (lut_lookup_not_36_nl));
      chn_lut_out_rsci_d_139_117 <= MUX1HOT_v_23_6_2(lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1,
          (lut_lookup_le_fraction_lpi_1_dfm_22[34:12]), (lut_lookup_le_fraction_lpi_1_dfm_9[34:12]),
          (lut_lookup_le_fraction_lpi_1_dfm_21[34:12]), (lut_lookup_lo_fraction_lpi_1_dfm_1[34:12]),
          (lut_lookup_lo_fraction_lpi_1_dfm_9[34:12]), {lut_lookup_lut_lookup_nor_16_cse
          , lut_lookup_and_29_cse , lut_lookup_and_30_cse , lut_lookup_and_31_cse
          , lut_lookup_and_132_cse , lut_lookup_and_133_cse});
      chn_lut_out_rsci_d_267_140 <= lut_in_data_sva_158;
      chn_lut_out_rsci_d_268 <= (lut_lookup_else_2_mux_1_nl) & (~ lut_lookup_1_and_svs_2);
      chn_lut_out_rsci_d_269 <= (lut_lookup_else_2_mux_27_nl) & (~ lut_lookup_2_and_svs_2);
      chn_lut_out_rsci_d_270 <= (lut_lookup_else_2_mux_53_nl) & (~ lut_lookup_3_and_svs_2);
      chn_lut_out_rsci_d_271 <= (lut_lookup_else_2_mux_79_nl) & (~ lut_lookup_4_and_svs_2);
      chn_lut_out_rsci_d_285_280 <= MUX1HOT_v_6_6_2(lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29,
          lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28, (lut_lookup_else_if_lut_lookup_else_if_and_2_nl),
          lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26, (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1[5:0]),
          (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13[5:0]), {lut_lookup_lut_lookup_nor_19_cse
          , lut_lookup_and_5_cse , lut_lookup_and_6_cse , lut_lookup_and_7_cse ,
          lut_lookup_and_138_cse , lut_lookup_and_139_cse});
      chn_lut_out_rsci_d_294_289 <= MUX1HOT_v_6_6_2(lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29,
          lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28, (lut_lookup_else_if_lut_lookup_else_if_and_5_nl),
          lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26, (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1[5:0]),
          (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13[5:0]), {lut_lookup_lut_lookup_nor_18_cse
          , lut_lookup_and_13_cse , lut_lookup_and_14_cse , lut_lookup_and_15_cse
          , lut_lookup_and_136_cse , lut_lookup_and_137_cse});
      chn_lut_out_rsci_d_303_298 <= MUX1HOT_v_6_6_2(lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29,
          lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28, (lut_lookup_else_if_lut_lookup_else_if_and_8_nl),
          lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26, (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1[5:0]),
          (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13[5:0]), {lut_lookup_lut_lookup_nor_17_cse
          , lut_lookup_and_21_cse , lut_lookup_and_22_cse , lut_lookup_and_23_cse
          , lut_lookup_and_134_cse , lut_lookup_and_135_cse});
      chn_lut_out_rsci_d_312_307 <= MUX1HOT_v_6_6_2(lut_lookup_le_index_0_5_0_lpi_1_dfm_29,
          lut_lookup_le_index_0_5_0_lpi_1_dfm_28, (lut_lookup_else_if_lut_lookup_else_if_and_11_nl),
          lut_lookup_le_index_0_5_0_lpi_1_dfm_26, (lut_lookup_lo_index_0_7_0_lpi_1_dfm_1[5:0]),
          (lut_lookup_lo_index_0_7_0_lpi_1_dfm_13[5:0]), {lut_lookup_lut_lookup_nor_16_cse
          , lut_lookup_and_29_cse , lut_lookup_and_30_cse , lut_lookup_and_31_cse
          , lut_lookup_and_132_cse , lut_lookup_and_133_cse});
      chn_lut_out_rsci_d_316 <= ~ lut_lookup_le_miss_1_sva;
      chn_lut_out_rsci_d_317 <= ~ lut_lookup_le_miss_2_sva;
      chn_lut_out_rsci_d_318 <= ~ lut_lookup_le_miss_3_sva;
      chn_lut_out_rsci_d_319 <= ~ lut_lookup_le_miss_sva;
      chn_lut_out_rsci_d_320 <= ~ lut_lookup_lo_miss_1_sva;
      chn_lut_out_rsci_d_321 <= ~ lut_lookup_lo_miss_2_sva;
      chn_lut_out_rsci_d_322 <= ~ lut_lookup_lo_miss_3_sva;
      chn_lut_out_rsci_d_323 <= ~ lut_lookup_lo_miss_sva;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_d_272 <= 1'b0;
      chn_lut_out_rsci_d_276 <= 1'b0;
      chn_lut_out_rsci_d_286 <= 1'b0;
      chn_lut_out_rsci_d_287 <= 1'b0;
      chn_lut_out_rsci_d_288 <= 1'b0;
    end
    else if ( chn_lut_out_and_13_cse ) begin
      chn_lut_out_rsci_d_272 <= MUX_s_1_2_2(lut_lookup_else_2_else_else_if_mux_5_itm_1,
          (lut_lookup_else_2_lut_lookup_else_2_and_4_nl), and_dcpl_59);
      chn_lut_out_rsci_d_276 <= MUX_s_1_2_2(cfg_lut_uflow_priority_1_sva_10, (lut_lookup_else_2_mux_103_nl),
          and_dcpl_59);
      chn_lut_out_rsci_d_286 <= MUX_s_1_2_2((lut_lookup_if_2_mux_21_nl), (lut_lookup_else_2_mux_107_nl),
          and_dcpl_59);
      chn_lut_out_rsci_d_287 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_8_nl),
          (lut_lookup_else_2_mux_108_nl), and_dcpl_59);
      chn_lut_out_rsci_d_288 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_9_nl),
          (lut_lookup_else_2_mux_109_nl), and_dcpl_59);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_d_273 <= 1'b0;
      chn_lut_out_rsci_d_277 <= 1'b0;
      chn_lut_out_rsci_d_295 <= 1'b0;
      chn_lut_out_rsci_d_296 <= 1'b0;
      chn_lut_out_rsci_d_297 <= 1'b0;
    end
    else if ( chn_lut_out_and_14_cse ) begin
      chn_lut_out_rsci_d_273 <= MUX_s_1_2_2(lut_lookup_else_2_else_else_if_mux_12_itm_1,
          (lut_lookup_else_2_lut_lookup_else_2_and_5_nl), and_dcpl_63);
      chn_lut_out_rsci_d_277 <= MUX_s_1_2_2(cfg_lut_uflow_priority_1_sva_10, (lut_lookup_else_2_mux_104_nl),
          and_dcpl_63);
      chn_lut_out_rsci_d_295 <= MUX_s_1_2_2((lut_lookup_if_2_mux_22_nl), (lut_lookup_else_2_mux_110_nl),
          and_dcpl_63);
      chn_lut_out_rsci_d_296 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_10_nl),
          (lut_lookup_else_2_mux_111_nl), and_dcpl_63);
      chn_lut_out_rsci_d_297 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_11_nl),
          (lut_lookup_else_2_mux_112_nl), and_dcpl_63);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_d_274 <= 1'b0;
      chn_lut_out_rsci_d_278 <= 1'b0;
      chn_lut_out_rsci_d_304 <= 1'b0;
      chn_lut_out_rsci_d_305 <= 1'b0;
      chn_lut_out_rsci_d_306 <= 1'b0;
    end
    else if ( chn_lut_out_and_15_cse ) begin
      chn_lut_out_rsci_d_274 <= MUX_s_1_2_2(lut_lookup_else_2_else_else_if_mux_19_itm_1,
          (lut_lookup_else_2_lut_lookup_else_2_and_6_nl), and_dcpl_67);
      chn_lut_out_rsci_d_278 <= MUX_s_1_2_2(cfg_lut_uflow_priority_1_sva_10, (lut_lookup_else_2_mux_105_nl),
          and_dcpl_67);
      chn_lut_out_rsci_d_304 <= MUX_s_1_2_2((lut_lookup_if_2_mux_23_nl), (lut_lookup_else_2_mux_113_nl),
          and_dcpl_67);
      chn_lut_out_rsci_d_305 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_12_nl),
          (lut_lookup_else_2_mux_114_nl), and_dcpl_67);
      chn_lut_out_rsci_d_306 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_13_nl),
          (lut_lookup_else_2_mux_115_nl), and_dcpl_67);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_lut_out_rsci_d_275 <= 1'b0;
      chn_lut_out_rsci_d_279 <= 1'b0;
      chn_lut_out_rsci_d_313 <= 1'b0;
      chn_lut_out_rsci_d_314 <= 1'b0;
      chn_lut_out_rsci_d_315 <= 1'b0;
    end
    else if ( chn_lut_out_and_16_cse ) begin
      chn_lut_out_rsci_d_275 <= MUX_s_1_2_2(lut_lookup_else_2_else_else_if_mux_26_itm_1,
          (lut_lookup_else_2_lut_lookup_else_2_and_7_nl), and_dcpl_71);
      chn_lut_out_rsci_d_279 <= MUX_s_1_2_2(cfg_lut_uflow_priority_1_sva_10, (lut_lookup_else_2_mux_106_nl),
          and_dcpl_71);
      chn_lut_out_rsci_d_313 <= MUX_s_1_2_2((lut_lookup_if_2_mux_24_nl), (lut_lookup_else_2_mux_116_nl),
          and_dcpl_71);
      chn_lut_out_rsci_d_314 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_14_nl),
          (lut_lookup_else_2_mux_117_nl), and_dcpl_71);
      chn_lut_out_rsci_d_315 <= MUX_s_1_2_2((lut_lookup_if_2_lut_lookup_if_2_and_15_nl),
          (lut_lookup_else_2_mux_118_nl), and_dcpl_71);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_lut_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_72 | and_dcpl_74) ) begin
      reg_chn_lut_out_rsci_ld_core_psct_cse <= ~ and_dcpl_74;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_1628 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_cfg_precision_1_sva_st_12_cse_1 <= 2'b0;
      reg_cfg_lut_le_function_1_sva_st_19_cse <= 1'b0;
      cfg_lut_le_index_offset_1_sva_4 <= 8'b0;
      cfg_lut_le_start_1_sva_41 <= 32'b0;
      lut_in_data_sva_154 <= 128'b0;
      cfg_lut_lo_start_1_sva_41 <= 32'b0;
      cfg_lut_le_index_select_1_sva_4 <= 8'b0;
      cfg_lut_lo_index_select_1_sva_4 <= 8'b0;
      lut_lookup_4_if_else_slc_32_svs_5 <= 1'b0;
      lut_lookup_3_if_else_slc_32_svs_5 <= 1'b0;
      lut_lookup_2_if_else_slc_32_svs_5 <= 1'b0;
      lut_lookup_1_if_else_slc_32_svs_5 <= 1'b0;
      cfg_lut_uflow_priority_1_sva_6 <= 1'b0;
      cfg_lut_oflow_priority_1_sva_6 <= 1'b0;
      cfg_lut_hybrid_priority_1_sva_6 <= 1'b0;
    end
    else if ( cfg_precision_and_cse ) begin
      reg_cfg_precision_1_sva_st_12_cse_1 <= cfg_precision_rsci_d;
      reg_cfg_lut_le_function_1_sva_st_19_cse <= cfg_lut_le_function_rsci_d;
      cfg_lut_le_index_offset_1_sva_4 <= cfg_lut_le_index_offset_rsci_d;
      cfg_lut_le_start_1_sva_41 <= cfg_lut_le_start_rsci_d;
      lut_in_data_sva_154 <= chn_lut_in_rsci_d_mxwt;
      cfg_lut_lo_start_1_sva_41 <= cfg_lut_lo_start_rsci_d;
      cfg_lut_le_index_select_1_sva_4 <= cfg_lut_le_index_select_rsci_d;
      cfg_lut_lo_index_select_1_sva_4 <= cfg_lut_lo_index_select_rsci_d;
      lut_lookup_4_if_else_slc_32_svs_5 <= lut_lookup_4_else_else_acc_1_itm_32;
      lut_lookup_3_if_else_slc_32_svs_5 <= lut_lookup_3_else_else_acc_1_itm_32;
      lut_lookup_2_if_else_slc_32_svs_5 <= lut_lookup_2_else_else_acc_1_itm_32;
      lut_lookup_1_if_else_slc_32_svs_5 <= lut_lookup_1_else_else_acc_1_itm_32;
      cfg_lut_uflow_priority_1_sva_6 <= cfg_lut_uflow_priority_rsci_d;
      cfg_lut_oflow_priority_1_sva_6 <= cfg_lut_oflow_priority_rsci_d;
      cfg_lut_hybrid_priority_1_sva_6 <= cfg_lut_hybrid_priority_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ mux_3_itm) ) begin
      reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[31]) ^ (cfg_lut_le_start_rsci_d[31]);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4 <= 8'b0;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 <= 1'b0;
      lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
      FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_2_is_addition_and_cse ) begin
      reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[31]) ^ (cfg_lut_lo_start_rsci_d[31]);
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[30:23]),
          (cfg_lut_lo_start_rsci_d[30:23]), and_dcpl_284);
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 <= IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0;
      lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
      FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3 <= readslicef_9_8_1((acc_6_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 <= 1'b0;
      reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse <= 1'b0;
      reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= 1'b0;
      FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_1_qr_lpi_1_dfm_5 <= 8'b0;
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 <= 1'b0;
      FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3 <= 8'b0;
      lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
      FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3 <= 8'b0;
      FpAdd_8U_23U_1_a_right_shift_qr_sva_3 <= 8'b0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_addition_and_1_cse ) begin
      reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[63]) ^ (cfg_lut_le_start_rsci_d[31]);
      reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[63]) ^ (cfg_lut_lo_start_rsci_d[31]);
      reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[95]) ^ (cfg_lut_le_start_rsci_d[31]);
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 <= ~(IsNaN_8U_23U_3_nor_10_tmp | (chn_lut_in_rsci_d_mxwt[94:87]!=8'b11111111));
      reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[95]) ^ (cfg_lut_lo_start_rsci_d[31]);
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse <= IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
      reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[127]) ^ (cfg_lut_le_start_rsci_d[31]);
      reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse
          <= (chn_lut_in_rsci_d_mxwt[127]) ^ (cfg_lut_lo_start_rsci_d[31]);
      FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[62:55]),
          (cfg_lut_le_start_rsci_d[30:23]), and_dcpl_288);
      FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[94:87]),
          (cfg_lut_le_start_rsci_d[30:23]), and_dcpl_296);
      FpAdd_8U_23U_1_qr_lpi_1_dfm_5 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[126:119]),
          (cfg_lut_le_start_rsci_d[30:23]), and_dcpl_304);
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 <= ~(IsNaN_8U_23U_3_nor_4_tmp | (chn_lut_in_rsci_d_mxwt[62:55]!=8'b11111111));
      FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3 <= readslicef_9_8_1((acc_8_nl));
      lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
      FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3 <= readslicef_9_8_1((acc_11_nl));
      FpAdd_8U_23U_1_a_right_shift_qr_sva_3 <= readslicef_9_8_1((acc_7_nl));
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 <= ~(IsNaN_8U_23U_8_nor_2_tmp_1 | IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & ((or_cse & main_stage_v_1) | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_lut_le_index_offset_1_sva_5 <= 8'b0;
      reg_cfg_precision_1_sva_st_13_cse_1 <= 2'b0;
      reg_cfg_lut_le_function_1_sva_st_20_cse <= 1'b0;
      cfg_lut_le_start_1_sva_2_30_0_1 <= 31'b0;
      cfg_lut_lo_start_1_sva_2_30_0_1 <= 31'b0;
      lut_in_data_sva_155 <= 128'b0;
      cfg_lut_le_index_select_1_sva_5 <= 8'b0;
      cfg_lut_lo_index_select_1_sva_5 <= 8'b0;
      lut_lookup_4_if_else_slc_32_svs_6 <= 1'b0;
      lut_lookup_3_if_else_slc_32_svs_6 <= 1'b0;
      lut_lookup_2_if_else_slc_32_svs_6 <= 1'b0;
      lut_lookup_1_if_else_slc_32_svs_6 <= 1'b0;
      cfg_lut_uflow_priority_1_sva_7 <= 1'b0;
      cfg_lut_oflow_priority_1_sva_7 <= 1'b0;
      cfg_lut_hybrid_priority_1_sva_7 <= 1'b0;
    end
    else if ( cfg_lut_le_index_offset_and_1_cse ) begin
      cfg_lut_le_index_offset_1_sva_5 <= cfg_lut_le_index_offset_1_sva_4;
      reg_cfg_precision_1_sva_st_13_cse_1 <= reg_cfg_precision_1_sva_st_12_cse_1;
      reg_cfg_lut_le_function_1_sva_st_20_cse <= reg_cfg_lut_le_function_1_sva_st_19_cse;
      cfg_lut_le_start_1_sva_2_30_0_1 <= cfg_lut_le_start_1_sva_41[30:0];
      cfg_lut_lo_start_1_sva_2_30_0_1 <= cfg_lut_lo_start_1_sva_41[30:0];
      lut_in_data_sva_155 <= lut_in_data_sva_154;
      cfg_lut_le_index_select_1_sva_5 <= cfg_lut_le_index_select_1_sva_4;
      cfg_lut_lo_index_select_1_sva_5 <= cfg_lut_lo_index_select_1_sva_4;
      lut_lookup_4_if_else_slc_32_svs_6 <= lut_lookup_4_if_else_slc_32_svs_5;
      lut_lookup_3_if_else_slc_32_svs_6 <= lut_lookup_3_if_else_slc_32_svs_5;
      lut_lookup_2_if_else_slc_32_svs_6 <= lut_lookup_2_if_else_slc_32_svs_5;
      lut_lookup_1_if_else_slc_32_svs_6 <= lut_lookup_1_if_else_slc_32_svs_5;
      cfg_lut_uflow_priority_1_sva_7 <= cfg_lut_uflow_priority_1_sva_6;
      cfg_lut_oflow_priority_1_sva_7 <= cfg_lut_oflow_priority_1_sva_6;
      cfg_lut_hybrid_priority_1_sva_7 <= cfg_lut_hybrid_priority_1_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm <= 2'b0;
    end
    else if ( and_dcpl_540 & (~ (reg_cfg_precision_1_sva_st_12_cse_1[0])) & or_cse
        & (reg_cfg_precision_1_sva_st_12_cse_1[1]) ) begin
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm <= FpAdd_8U_23U_1_mux1h_1_itm[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm <= 6'b0;
    end
    else if ( (and_956_cse | (FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 & (~
        reg_cfg_lut_le_function_1_sva_st_19_cse))) & and_dcpl_540 & or_cse ) begin
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm <= FpAdd_8U_23U_1_mux1h_1_itm[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_1_sva_3 <= 50'b0;
    end
    else if ( core_wen & (and_284_rgt | and_286_rgt | and_288_rgt | and_290_rgt)
        & not_tmp_47 ) begin
      FpAdd_8U_23U_1_int_mant_p1_1_sva_3 <= MUX1HOT_v_50_4_2((lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl),
          (lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl), (lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl),
          (lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl), {and_284_rgt , and_286_rgt , and_288_rgt
          , and_290_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 <= 8'b0;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_2_and_35_cse ) begin
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 <= FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 <= IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
      IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 <= IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_int_mant_p1_1_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_cse & (~ reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse))
        | and_292_rgt) & (~ mux_20_itm) ) begin
      FpAdd_8U_23U_2_int_mant_p1_1_sva_3 <= MUX_v_50_2_2((lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl),
          (lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl), and_292_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm <= 2'b0;
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm <= 2'b0;
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm <= 2'b0;
    end
    else if ( and_961_cse ) begin
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm <= FpAdd_8U_23U_1_mux1h_3_itm[7:6];
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm <= FpAdd_8U_23U_1_mux1h_5_itm[7:6];
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm <= FpAdd_8U_23U_1_mux1h_7_itm[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm <= 6'b0;
    end
    else if ( (and_956_cse | (FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 & (~
        reg_cfg_lut_le_function_1_sva_st_19_cse))) & and_dcpl_540 & or_cse ) begin
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm <= FpAdd_8U_23U_1_mux1h_3_itm[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_2_sva_3 <= 50'b0;
    end
    else if ( core_wen & (and_300_rgt | and_302_rgt | and_304_rgt | and_306_rgt)
        & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_1_int_mant_p1_2_sva_3 <= MUX1HOT_v_50_4_2((lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl),
          (lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl), (lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl),
          (lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl), {and_300_rgt , and_302_rgt , and_304_rgt
          , and_306_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 <= 8'b0;
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_2_and_36_cse ) begin
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 <= FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4;
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 <= IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_int_mant_p1_2_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_cse & (~ reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse))
        | and_308_rgt) & (~ mux_26_itm) ) begin
      FpAdd_8U_23U_2_int_mant_p1_2_sva_3 <= MUX_v_50_2_2((lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl),
          (lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl), and_308_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm <= 6'b0;
    end
    else if ( (and_956_cse | ((~ reg_cfg_lut_le_function_1_sva_st_19_cse) & FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5))
        & and_dcpl_540 & or_cse ) begin
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm <= FpAdd_8U_23U_1_mux1h_5_itm[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_3_sva_3 <= 50'b0;
    end
    else if ( core_wen & (and_316_rgt | and_318_rgt | and_320_rgt | and_322_rgt)
        & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_1_int_mant_p1_3_sva_3 <= MUX1HOT_v_50_4_2((lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl),
          (lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl), (lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl),
          (lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl), {and_316_rgt , and_318_rgt , and_320_rgt
          , and_322_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 <= 8'b0;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 <= 1'b0;
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse <= 1'b0;
      FpAdd_8U_23U_2_qr_lpi_1_dfm_5 <= 8'b0;
      IsNaN_8U_23U_8_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_2_and_37_cse ) begin
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 <= FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 <= IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse <= reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
      FpAdd_8U_23U_2_qr_lpi_1_dfm_5 <= FpAdd_8U_23U_2_qr_lpi_1_dfm_4;
      IsNaN_8U_23U_8_land_lpi_1_dfm_4 <= nor_469_cse;
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 <= nor_482_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_int_mant_p1_3_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_cse & (~ reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse))
        | and_324_rgt) & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_2_int_mant_p1_3_sva_3 <= MUX_v_50_2_2((lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl),
          (lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl), and_324_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm <= 6'b0;
    end
    else if ( (and_956_cse | ((~ reg_cfg_lut_le_function_1_sva_st_19_cse) & FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5))
        & and_dcpl_540 & or_cse ) begin
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm <= FpAdd_8U_23U_1_mux1h_7_itm[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_sva_3 <= 50'b0;
    end
    else if ( core_wen & (and_330_rgt | and_332_rgt | and_334_rgt | and_336_rgt)
        & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_1_int_mant_p1_sva_3 <= MUX1HOT_v_50_4_2((lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl),
          (lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl), (lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl),
          (lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl), {and_330_rgt , and_332_rgt , and_334_rgt
          , and_336_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_int_mant_p1_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_cse & (~ reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse))
        | and_338_rgt) & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_2_int_mant_p1_sva_3 <= MUX_v_50_2_2((lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl),
          (lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl), and_338_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & ((or_cse & main_stage_v_2) | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_lut_le_start_1_sva_3_30_0_1 <= 31'b0;
      lut_in_data_sva_156 <= 128'b0;
      cfg_precision_1_sva_st_70 <= 2'b0;
      cfg_lut_le_function_1_sva_st_41 <= 1'b0;
      cfg_lut_le_index_offset_1_sva_6 <= 8'b0;
      cfg_lut_le_index_select_1_sva_6 <= 8'b0;
      cfg_lut_lo_index_select_1_sva_6 <= 8'b0;
      lut_lookup_if_else_else_slc_10_mdf_1_sva_3 <= 1'b0;
      lut_lookup_1_if_else_slc_32_svs_7 <= 1'b0;
      lut_lookup_if_else_else_slc_10_mdf_2_sva_3 <= 1'b0;
      lut_lookup_2_if_else_slc_32_svs_7 <= 1'b0;
      lut_lookup_if_else_else_slc_10_mdf_3_sva_3 <= 1'b0;
      lut_lookup_3_if_else_slc_32_svs_7 <= 1'b0;
      lut_lookup_if_else_else_slc_10_mdf_sva_3 <= 1'b0;
      lut_lookup_4_if_else_slc_32_svs_7 <= 1'b0;
      cfg_lut_uflow_priority_1_sva_8 <= 1'b0;
      cfg_lut_oflow_priority_1_sva_8 <= 1'b0;
      cfg_lut_hybrid_priority_1_sva_8 <= 1'b0;
    end
    else if ( cfg_lut_le_start_and_cse ) begin
      cfg_lut_le_start_1_sva_3_30_0_1 <= cfg_lut_le_start_1_sva_2_30_0_1;
      lut_in_data_sva_156 <= lut_in_data_sva_155;
      cfg_precision_1_sva_st_70 <= reg_cfg_precision_1_sva_st_13_cse_1;
      cfg_lut_le_function_1_sva_st_41 <= reg_cfg_lut_le_function_1_sva_st_20_cse;
      cfg_lut_le_index_offset_1_sva_6 <= cfg_lut_le_index_offset_1_sva_5;
      cfg_lut_le_index_select_1_sva_6 <= cfg_lut_le_index_select_1_sva_5;
      cfg_lut_lo_index_select_1_sva_6 <= cfg_lut_lo_index_select_1_sva_5;
      lut_lookup_if_else_else_slc_10_mdf_1_sva_3 <= lut_lookup_1_if_else_else_acc_itm_10;
      lut_lookup_1_if_else_slc_32_svs_7 <= lut_lookup_1_if_else_slc_32_svs_6;
      lut_lookup_if_else_else_slc_10_mdf_2_sva_3 <= lut_lookup_2_if_else_else_acc_itm_10;
      lut_lookup_2_if_else_slc_32_svs_7 <= lut_lookup_2_if_else_slc_32_svs_6;
      lut_lookup_if_else_else_slc_10_mdf_3_sva_3 <= lut_lookup_3_if_else_else_acc_itm_10;
      lut_lookup_3_if_else_slc_32_svs_7 <= lut_lookup_3_if_else_slc_32_svs_6;
      lut_lookup_if_else_else_slc_10_mdf_sva_3 <= lut_lookup_4_if_else_else_acc_itm_10;
      lut_lookup_4_if_else_slc_32_svs_7 <= lut_lookup_4_if_else_slc_32_svs_6;
      cfg_lut_uflow_priority_1_sva_8 <= cfg_lut_uflow_priority_1_sva_7;
      cfg_lut_oflow_priority_1_sva_8 <= cfg_lut_oflow_priority_1_sva_7;
      cfg_lut_hybrid_priority_1_sva_8 <= cfg_lut_hybrid_priority_1_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (and_344_rgt | and_dcpl_148 | and_347_rgt) & (~ (mux_39_nl))
        ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_1_lpi_1_dfm_4, lut_lookup_1_if_else_else_acc_itm_10,
          {and_344_rgt , and_dcpl_148 , and_347_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= 1'b0;
    end
    else if ( (~ (mux_1219_nl)) & core_wen ) begin
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= lut_lookup_if_else_else_else_le_index_s_1_sva[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= 2'b0;
    end
    else if ( or_66_cse & IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & or_cse & (~(lut_lookup_1_if_else_else_acc_itm_10
        | reg_cfg_lut_le_function_1_sva_st_20_cse)) & and_dcpl_576 ) begin
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= lut_lookup_if_else_else_else_le_index_s_1_sva[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= 23'b0;
      FpMantRNE_49U_24U_1_else_carry_1_sva_2 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_o_mant_and_cse ) begin
      lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[47:25];
      FpMantRNE_49U_24U_1_else_carry_1_sva_2 <= FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm <= 2'b0;
    end
    else if ( or_1936_cse & and_dcpl_576 & (reg_cfg_precision_1_sva_st_13_cse_1[1])
        & nor_865_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm <= MUX1HOT_v_2_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl),
          reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm, (lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt[7:6]),
          {FpAdd_8U_23U_o_expo_and_3_ssc , FpAdd_8U_23U_and_51_ssc , FpAdd_8U_23U_and_43_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm <= 6'b0;
    end
    else if ( (~ (mux_1224_nl)) & and_dcpl_576 & or_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm <= MUX1HOT_v_6_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl),
          reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm, (lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt[5:0]),
          {FpAdd_8U_23U_o_expo_and_3_ssc , (FpAdd_8U_23U_o_expo_or_3_nl) , FpAdd_8U_23U_and_43_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_13_itm_4 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse & (mux_59_nl) ) begin
      FpAdd_8U_23U_1_mux_13_itm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_13_itm_3, lut_lookup_1_else_else_else_if_acc_itm_3_1,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6 <= 1'b0;
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6 <= 1'b0;
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6 <= 1'b0;
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_3_land_lpi_1_dfm_st_6 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_6_cse ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7,
          IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5, and_dcpl_162);
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6 <= MUX_s_1_2_2(IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5,
          IsNaN_8U_23U_4_land_1_lpi_1_dfm_4, and_dcpl_162);
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_7,
          IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5, and_dcpl_162);
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6 <= MUX_s_1_2_2(IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5,
          IsNaN_8U_23U_4_land_2_lpi_1_dfm_5, and_dcpl_162);
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7,
          IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5, and_dcpl_162);
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6 <= MUX_s_1_2_2(IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5,
          IsNaN_8U_23U_4_land_3_lpi_1_dfm_5, and_dcpl_162);
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_lpi_1_dfm_7,
          reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse, and_dcpl_162);
      IsNaN_8U_23U_3_land_lpi_1_dfm_st_6 <= MUX_s_1_2_2(reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse,
          IsNaN_8U_23U_4_land_lpi_1_dfm_4, and_dcpl_162);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
      IsNaN_8U_23U_8_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 <= 1'b0;
      lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
      reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
      reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 <= 1'b0;
      lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
      reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
      IsNaN_8U_23U_8_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_8U_23U_7_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_lpi_1_dfm_st_6 <= 1'b0;
      lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_and_cse ) begin
      reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
      IsNaN_8U_23U_8_land_1_lpi_1_dfm_7 <= IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 <= IsNaN_8U_23U_7_land_1_lpi_1_dfm_6;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 <= IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
      lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2 <= lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp;
      reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp;
      reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp;
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 <= IsNaN_8U_23U_8_land_3_lpi_1_dfm_4;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 <= IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 <= IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
      lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2 <= lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp;
      reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp;
      IsNaN_8U_23U_8_land_lpi_1_dfm_5 <= IsNaN_8U_23U_8_land_lpi_1_dfm_4;
      IsNaN_8U_23U_7_land_lpi_1_dfm_7 <= IsNaN_8U_23U_7_land_lpi_1_dfm_6;
      IsNaN_8U_23U_7_land_lpi_1_dfm_st_6 <= reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
      lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2 <= lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse & mux_tmp_35 ) begin
      FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 <= MUX_s_1_2_2(nor_5_cse_1, IsNaN_8U_23U_1_land_1_lpi_1_dfm_7,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_61_nl) ) begin
      lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[47:25];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_49U_24U_2_else_carry_1_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_66_nl) ) begin
      FpMantRNE_49U_24U_2_else_carry_1_sva_2 <= MUX_s_1_2_2(FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0,
          (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12 <= 8'b0;
    end
    else if ( core_wen & (FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt | FpAdd_8U_23U_2_and_4_rgt
        | FpAdd_8U_23U_2_and_5_rgt) & (~ (mux_69_nl)) ) begin
      FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12 <= MUX1HOT_v_8_3_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_nl),
          FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5, (lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl),
          {FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt , FpAdd_8U_23U_2_and_4_rgt
          , FpAdd_8U_23U_2_and_5_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_lut_lo_start_1_sva_3_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_82_nl)) ) begin
      cfg_lut_lo_start_1_sva_3_30_0_1 <= cfg_lut_lo_start_1_sva_2_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_13_itm_3 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_86_nl) ) begin
      FpAdd_8U_23U_2_mux_13_itm_3 <= MUX_s_1_2_2(FpAdd_8U_23U_2_mux_13_itm_1, (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_2_is_inf_and_cse ) begin
      FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 <= MUX_s_1_2_2(nor_13_cse, IsNaN_8U_23U_7_land_1_lpi_1_dfm_6,
          and_dcpl_161);
      FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 <= MUX_s_1_2_2(nor_31_cse, IsNaN_8U_23U_7_land_2_lpi_1_dfm_6,
          and_dcpl_161);
      FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 <= MUX_s_1_2_2(nor_42_cse, IsNaN_8U_23U_7_land_3_lpi_1_dfm_6,
          and_dcpl_161);
      FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 <= MUX_s_1_2_2(nor_54_cse, IsNaN_8U_23U_7_land_lpi_1_dfm_6,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse & (~
        (mux_89_nl)) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_2_lpi_1_dfm_5, lut_lookup_2_if_else_else_acc_itm_10,
          {and_364_rgt , and_dcpl_148 , and_347_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= 1'b0;
    end
    else if ( (~ (mux_1226_nl)) & core_wen ) begin
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= lut_lookup_if_else_else_else_le_index_s_2_sva[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= 2'b0;
    end
    else if ( or_66_cse & IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & or_cse & (~(lut_lookup_2_if_else_else_acc_itm_10
        | reg_cfg_lut_le_function_1_sva_st_20_cse)) & and_dcpl_576 ) begin
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= lut_lookup_if_else_else_else_le_index_s_2_sva[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= 23'b0;
      FpMantRNE_49U_24U_1_else_carry_2_sva_2 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_o_mant_and_1_cse ) begin
      lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[47:25];
      FpMantRNE_49U_24U_1_else_carry_2_sva_2 <= FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm <= 2'b0;
    end
    else if ( (nor_855_cse | lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp) & and_dcpl_576
        & (reg_cfg_precision_1_sva_st_13_cse_1[1]) & nor_865_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm <= MUX1HOT_v_2_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl),
          reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm, (lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt[7:6]),
          {FpAdd_8U_23U_o_expo_and_2_ssc , FpAdd_8U_23U_and_53_ssc , FpAdd_8U_23U_and_45_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm <= 6'b0;
    end
    else if ( (~ (mux_1230_nl)) & and_dcpl_576 & or_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm <= MUX1HOT_v_6_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_10_nl),
          reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm, (lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt[5:0]),
          {FpAdd_8U_23U_o_expo_and_2_ssc , (FpAdd_8U_23U_o_expo_or_2_nl) , FpAdd_8U_23U_and_45_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_29_itm_4 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse & (mux_121_nl) )
        begin
      FpAdd_8U_23U_1_mux_29_itm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_29_itm_3, lut_lookup_2_else_else_else_if_acc_itm_3_1,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 <= 1'b0;
      FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 <= 1'b0;
      FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_inf_and_1_cse ) begin
      FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 <= MUX_s_1_2_2(nor_27_cse_1, IsNaN_8U_23U_1_land_2_lpi_1_dfm_7,
          and_dcpl_161);
      FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 <= MUX_s_1_2_2(nor_38_cse_1, IsNaN_8U_23U_1_land_3_lpi_1_dfm_7,
          and_dcpl_161);
      FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 <= MUX_s_1_2_2(nor_50_cse_1, IsNaN_8U_23U_1_land_lpi_1_dfm_7,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_123_nl) ) begin
      lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[47:25];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_49U_24U_2_else_carry_2_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_128_nl) ) begin
      FpMantRNE_49U_24U_2_else_carry_2_sva_2 <= MUX_s_1_2_2(FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0,
          (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12 <= 8'b0;
    end
    else if ( core_wen & (FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt |
        FpAdd_8U_23U_2_and_10_rgt | FpAdd_8U_23U_2_and_11_rgt) & (~ (mux_131_nl))
        ) begin
      FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12 <= MUX1HOT_v_8_3_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_2_nl),
          FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5, (lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl),
          {FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt , FpAdd_8U_23U_2_and_10_rgt
          , FpAdd_8U_23U_2_and_11_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6 <= 1'b0;
      lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_8_aelse_and_1_cse ) begin
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 <= IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 <= IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6 <= IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
      lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2 <= lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_29_itm_3 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_135_nl) ) begin
      FpAdd_8U_23U_2_mux_29_itm_3 <= MUX_s_1_2_2(FpAdd_8U_23U_2_mux_29_itm_1, (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse & (~
        (mux_138_nl)) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_3_lpi_1_dfm_5, lut_lookup_3_if_else_else_acc_itm_10,
          {and_364_rgt , and_dcpl_148 , and_347_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= 1'b0;
    end
    else if ( (~ (mux_1232_nl)) & core_wen ) begin
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= lut_lookup_if_else_else_else_le_index_s_3_sva[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= 2'b0;
    end
    else if ( or_66_cse & IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & or_cse & (~(lut_lookup_3_if_else_else_acc_itm_10
        | reg_cfg_lut_le_function_1_sva_st_20_cse)) & and_dcpl_576 ) begin
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= lut_lookup_if_else_else_else_le_index_s_3_sva[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= 23'b0;
      FpMantRNE_49U_24U_1_else_carry_3_sva_2 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_o_mant_and_2_cse ) begin
      lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[47:25];
      FpMantRNE_49U_24U_1_else_carry_3_sva_2 <= FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm <= 2'b0;
    end
    else if ( ((~((mux_1233_nl) | nor_38_cse_1 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_7))
        | lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp) & and_dcpl_576 & (reg_cfg_precision_1_sva_st_13_cse_1[1])
        & nor_865_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm <= MUX1HOT_v_2_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl),
          reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm, (lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt[7:6]),
          {FpAdd_8U_23U_o_expo_and_1_ssc , FpAdd_8U_23U_and_55_ssc , FpAdd_8U_23U_and_47_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm <= 6'b0;
    end
    else if ( (~ (mux_1237_nl)) & and_dcpl_576 & or_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm <= MUX1HOT_v_6_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl),
          reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm, (lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt[5:0]),
          {FpAdd_8U_23U_o_expo_and_1_ssc , (FpAdd_8U_23U_o_expo_or_1_nl) , FpAdd_8U_23U_and_47_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_45_itm_4 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse & (mux_157_nl) )
        begin
      FpAdd_8U_23U_1_mux_45_itm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_45_itm_3, lut_lookup_3_else_else_else_if_acc_itm_3_1,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_159_nl) ) begin
      lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[47:25];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_49U_24U_2_else_carry_3_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_164_nl) ) begin
      FpMantRNE_49U_24U_2_else_carry_3_sva_2 <= MUX_s_1_2_2(FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0,
          (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12 <= 8'b0;
    end
    else if ( core_wen & (FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt |
        FpAdd_8U_23U_2_and_16_rgt | FpAdd_8U_23U_2_and_17_rgt) & (~ (mux_167_nl))
        ) begin
      FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12 <= MUX1HOT_v_8_3_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_4_nl),
          FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5, (lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl),
          {FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt , FpAdd_8U_23U_2_and_16_rgt
          , FpAdd_8U_23U_2_and_17_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_45_itm_3 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_171_nl) ) begin
      FpAdd_8U_23U_2_mux_45_itm_3 <= MUX_s_1_2_2(FpAdd_8U_23U_2_mux_45_itm_1, (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse & (~
        (mux_174_nl)) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_1_land_lpi_1_dfm_7,
          IsNaN_8U_23U_4_land_lpi_1_dfm_4, lut_lookup_4_if_else_else_acc_itm_10,
          {and_364_rgt , and_dcpl_148 , and_347_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= 1'b0;
    end
    else if ( (~ (mux_1239_nl)) & core_wen ) begin
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm
          <= lut_lookup_if_else_else_else_le_index_s_sva[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= 2'b0;
    end
    else if ( or_66_cse & IsNaN_8U_23U_1_land_lpi_1_dfm_7 & or_cse & (~(lut_lookup_4_if_else_else_acc_itm_10
        | reg_cfg_lut_le_function_1_sva_st_20_cse)) & and_dcpl_576 ) begin
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm
          <= lut_lookup_if_else_else_else_le_index_s_sva[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= 23'b0;
      FpMantRNE_49U_24U_1_else_carry_sva_2 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_o_mant_and_3_cse ) begin
      lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2
          <= FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[47:25];
      FpMantRNE_49U_24U_1_else_carry_sva_2 <= FpMantRNE_49U_24U_1_else_carry_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm <= 2'b0;
    end
    else if ( ((~((mux_1240_nl) | nor_50_cse_1 | IsNaN_8U_23U_1_land_lpi_1_dfm_7))
        | lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp) & and_dcpl_576 & (reg_cfg_precision_1_sva_st_13_cse_1[1])
        & nor_865_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm <= MUX1HOT_v_2_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl),
          reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm, (lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt[7:6]),
          {FpAdd_8U_23U_o_expo_and_ssc , FpAdd_8U_23U_and_57_ssc , FpAdd_8U_23U_and_49_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm <= 6'b0;
    end
    else if ( (~ (mux_1244_nl)) & and_dcpl_576 & or_cse ) begin
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm <= MUX1HOT_v_6_3_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_8_nl),
          reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm, (lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt[5:0]),
          {FpAdd_8U_23U_o_expo_and_ssc , (FpAdd_8U_23U_o_expo_or_nl) , FpAdd_8U_23U_and_49_ssc});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_61_itm_4 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse & (mux_200_nl) )
        begin
      FpAdd_8U_23U_1_mux_61_itm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_61_itm_3, lut_lookup_4_else_else_else_if_acc_itm_3_1,
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_202_nl) ) begin
      lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2
          <= FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[47:25];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_49U_24U_2_else_carry_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_207_nl) ) begin
      FpMantRNE_49U_24U_2_else_carry_sva_2 <= MUX_s_1_2_2(FpMantRNE_49U_24U_2_else_carry_sva_mx0w0,
          (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12 <= 8'b0;
    end
    else if ( core_wen & (FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt |
        FpAdd_8U_23U_2_and_22_rgt | FpAdd_8U_23U_2_and_23_rgt) & (~ (mux_211_nl))
        ) begin
      FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12 <= MUX1HOT_v_8_3_2((FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_6_nl),
          FpAdd_8U_23U_2_qr_lpi_1_dfm_5, (lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl),
          {FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt , FpAdd_8U_23U_2_and_22_rgt
          , FpAdd_8U_23U_2_and_23_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_61_itm_3 <= 1'b0;
    end
    else if ( core_wen & FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse
        & (mux_215_nl) ) begin
      FpAdd_8U_23U_2_mux_61_itm_3 <= MUX_s_1_2_2(FpAdd_8U_23U_2_mux_61_itm_1, (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8]),
          and_dcpl_161);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & ((or_cse & main_stage_v_3) | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_lut_le_index_offset_1_sva_7 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) ) begin
      cfg_lut_le_index_offset_1_sva_7 <= cfg_lut_le_index_offset_1_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse
        & (~ (mux_218_nl)) ) begin
      lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= MUX_s_1_2_2(lut_lookup_1_if_else_else_else_else_acc_itm_32_1, lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1,
          and_428_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_219_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_if_else_slc_32_svs_st_5 <= 1'b0;
      lut_lookup_2_if_else_slc_32_svs_st_5 <= 1'b0;
      lut_lookup_3_if_else_slc_32_svs_st_5 <= 1'b0;
      lut_lookup_4_if_else_slc_32_svs_st_5 <= 1'b0;
    end
    else if ( lut_lookup_if_else_if_and_cse ) begin
      lut_lookup_1_if_else_slc_32_svs_st_5 <= FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
      lut_lookup_2_if_else_slc_32_svs_st_5 <= FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
      lut_lookup_3_if_else_slc_32_svs_st_5 <= FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
      lut_lookup_4_if_else_slc_32_svs_st_5 <= FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_71 <= 2'b0;
      cfg_lut_le_function_1_sva_st_42 <= 1'b0;
      cfg_lut_hybrid_priority_1_sva_9 <= 1'b0;
      cfg_lut_uflow_priority_1_sva_9 <= 1'b0;
      lut_lookup_else_unequal_tmp_18 <= 1'b0;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_25 <= 6'b0;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_27 <= 6'b0;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25 <= 6'b0;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27 <= 6'b0;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25 <= 6'b0;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27 <= 6'b0;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25 <= 6'b0;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27 <= 6'b0;
      cfg_lut_oflow_priority_1_sva_9 <= 1'b0;
      lut_in_data_sva_157 <= 128'b0;
    end
    else if ( cfg_precision_and_24_cse ) begin
      cfg_precision_1_sva_st_71 <= cfg_precision_1_sva_st_70;
      cfg_lut_le_function_1_sva_st_42 <= cfg_lut_le_function_1_sva_st_41;
      cfg_lut_hybrid_priority_1_sva_9 <= cfg_lut_hybrid_priority_1_sva_8;
      cfg_lut_uflow_priority_1_sva_9 <= cfg_lut_uflow_priority_1_sva_8;
      lut_lookup_else_unequal_tmp_18 <= lut_lookup_unequal_tmp_mx0w0;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_25 <= MUX_v_6_2_2(6'b000000, lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2,
          lut_lookup_else_else_slc_32_mdf_sva_7);
      lut_lookup_le_index_0_5_0_lpi_1_dfm_27 <= lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          & ({{5{lut_lookup_4_if_else_else_else_if_acc_itm_3_1}}, lut_lookup_4_if_else_else_else_if_acc_itm_3_1})
          & (signext_6_1(~ lut_lookup_if_else_else_slc_10_mdf_sva_3)) & ({{5{lut_lookup_4_if_else_slc_32_svs_7}},
          lut_lookup_4_if_else_slc_32_svs_7});
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25 <= MUX_v_6_2_2(6'b000000, lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2,
          lut_lookup_else_else_slc_32_mdf_3_sva_7);
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27 <= lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          & ({{5{lut_lookup_3_if_else_else_else_if_acc_itm_3_1}}, lut_lookup_3_if_else_else_else_if_acc_itm_3_1})
          & (signext_6_1(~ lut_lookup_if_else_else_slc_10_mdf_3_sva_3)) & ({{5{lut_lookup_3_if_else_slc_32_svs_7}},
          lut_lookup_3_if_else_slc_32_svs_7});
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25 <= MUX_v_6_2_2(6'b000000, lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2,
          lut_lookup_else_else_slc_32_mdf_2_sva_7);
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27 <= lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          & ({{5{lut_lookup_2_if_else_else_else_if_acc_itm_3_1}}, lut_lookup_2_if_else_else_else_if_acc_itm_3_1})
          & (signext_6_1(~ lut_lookup_if_else_else_slc_10_mdf_2_sva_3)) & ({{5{lut_lookup_2_if_else_slc_32_svs_7}},
          lut_lookup_2_if_else_slc_32_svs_7});
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25 <= MUX_v_6_2_2(6'b000000, lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2,
          lut_lookup_else_else_slc_32_mdf_1_sva_7);
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27 <= lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          & ({{5{lut_lookup_1_if_else_else_else_if_acc_itm_3}}, lut_lookup_1_if_else_else_else_if_acc_itm_3})
          & (signext_6_1(~ lut_lookup_if_else_else_slc_10_mdf_1_sva_3)) & ({{5{lut_lookup_1_if_else_slc_32_svs_7}},
          lut_lookup_1_if_else_slc_32_svs_7});
      cfg_lut_oflow_priority_1_sva_9 <= cfg_lut_oflow_priority_1_sva_8;
      lut_in_data_sva_157 <= lut_in_data_sva_156;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1 <= 1'b0;
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1 <= ~ (cfg_lut_le_index_select_1_sva_6[0]);
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= z_out_4[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_1_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse & (mux_225_nl)
        ) begin
      lut_lookup_else_else_else_asn_mdf_1_sva_st_3 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_13_itm_4,
          lut_lookup_1_if_else_else_else_if_acc_itm_3, and_430_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1 <= 1'b0;
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1 <= ~ (cfg_lut_lo_index_select_1_sva_6[0]);
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_228_nl) ) begin
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= FpAdd_8U_23U_2_mux_13_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse
        & (~ (mux_231_nl)) ) begin
      lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= MUX_s_1_2_2(lut_lookup_2_if_else_else_else_else_acc_itm_32_1, lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1,
          and_428_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_232_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1 <= 1'b0;
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1 <= ~ (cfg_lut_le_index_select_1_sva_6[0]);
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= z_out_5[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_2_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse & (mux_237_nl)
        ) begin
      lut_lookup_else_else_else_asn_mdf_2_sva_st_3 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_29_itm_4,
          lut_lookup_2_if_else_else_else_if_acc_itm_3_1, and_430_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1 <= 1'b0;
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1 <= ~ (cfg_lut_lo_index_select_1_sva_6[0]);
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_240_nl) ) begin
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= FpAdd_8U_23U_2_mux_29_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse
        & (~ (mux_244_nl)) ) begin
      lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= MUX_s_1_2_2(lut_lookup_3_if_else_else_else_else_acc_itm_32_1, lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1,
          and_428_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_245_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1 <= 1'b0;
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1 <= ~ (cfg_lut_le_index_select_1_sva_6[0]);
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= z_out_6[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_3_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse & (mux_250_nl)
        ) begin
      lut_lookup_else_else_else_asn_mdf_3_sva_st_3 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_45_itm_4,
          lut_lookup_3_if_else_else_else_if_acc_itm_3_1, and_430_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1 <= 1'b0;
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1 <= ~ (cfg_lut_lo_index_select_1_sva_6[0]);
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_253_nl) ) begin
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= FpAdd_8U_23U_2_mux_45_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse
        & (~ (mux_256_nl)) ) begin
      lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
          <= MUX_s_1_2_2(lut_lookup_4_if_else_else_else_else_acc_itm_32_1, lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1,
          and_428_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_257_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_sva_st_3 <= IsNaN_8U_23U_1_land_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1 <= 1'b0;
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1 <= ~ (cfg_lut_le_index_select_1_sva_6[0]);
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= z_out_7[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_sva_st_3 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse & (mux_262_nl)
        ) begin
      lut_lookup_else_else_else_asn_mdf_sva_st_3 <= MUX_s_1_2_2(FpAdd_8U_23U_1_mux_61_itm_4,
          lut_lookup_4_if_else_else_else_if_acc_itm_3_1, and_430_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1 <= 1'b0;
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b0;
    end
    else if ( FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1 <= ~ (cfg_lut_lo_index_select_1_sva_6[0]);
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_265_nl) ) begin
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
          <= FpAdd_8U_23U_2_mux_61_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_5 <= 1'b0;
    end
    else if ( core_wen & ((or_cse & main_stage_v_4) | main_stage_v_5_mx0c1) ) begin
      main_stage_v_5 <= ~ main_stage_v_5_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_lut_hybrid_priority_1_sva_10 <= 1'b0;
      cfg_lut_oflow_priority_1_sva_10 <= 1'b0;
      lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1 <= 23'b0;
      lut_lookup_le_fraction_1_lpi_1_dfm_22 <= 35'b0;
      lut_lookup_le_fraction_1_lpi_1_dfm_21 <= 35'b0;
      lut_lookup_lo_fraction_1_lpi_1_dfm_9 <= 35'b0;
      lut_lookup_unequal_tmp_13 <= 1'b0;
      lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1 <= 23'b0;
      lut_lookup_le_fraction_2_lpi_1_dfm_22 <= 35'b0;
      lut_lookup_le_fraction_2_lpi_1_dfm_21 <= 35'b0;
      lut_lookup_lo_fraction_2_lpi_1_dfm_9 <= 35'b0;
      lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1 <= 23'b0;
      lut_lookup_le_fraction_3_lpi_1_dfm_22 <= 35'b0;
      lut_lookup_le_fraction_3_lpi_1_dfm_21 <= 35'b0;
      lut_lookup_lo_fraction_3_lpi_1_dfm_9 <= 35'b0;
      lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1 <= 23'b0;
      lut_lookup_le_fraction_lpi_1_dfm_22 <= 35'b0;
      lut_lookup_le_fraction_lpi_1_dfm_21 <= 35'b0;
      lut_lookup_lo_fraction_lpi_1_dfm_9 <= 35'b0;
      lut_in_data_sva_158 <= 128'b0;
      lut_lookup_1_and_svs_2 <= 1'b0;
      lut_lookup_2_and_svs_2 <= 1'b0;
      lut_lookup_3_and_svs_2 <= 1'b0;
      cfg_lut_uflow_priority_1_sva_10 <= 1'b0;
      lut_lookup_4_and_svs_2 <= 1'b0;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_29 <= 6'b0;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_28 <= 6'b0;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_26 <= 6'b0;
      lut_lookup_else_unequal_tmp_13 <= 1'b0;
      cfg_lut_le_function_1_sva_10 <= 1'b0;
      reg_lut_lookup_if_unequal_cse <= 1'b0;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29 <= 6'b0;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28 <= 6'b0;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26 <= 6'b0;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29 <= 6'b0;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28 <= 6'b0;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26 <= 6'b0;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29 <= 6'b0;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28 <= 6'b0;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26 <= 6'b0;
      lut_lookup_lo_uflow_lpi_1_dfm_4 <= 1'b0;
      cfg_precision_1_sva_st_107 <= 2'b0;
      lut_lookup_lo_uflow_3_lpi_1_dfm_4 <= 1'b0;
      lut_lookup_lo_uflow_2_lpi_1_dfm_4 <= 1'b0;
      lut_lookup_lo_uflow_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( cfg_lut_hybrid_priority_and_cse ) begin
      cfg_lut_hybrid_priority_1_sva_10 <= cfg_lut_hybrid_priority_1_sva_9;
      cfg_lut_oflow_priority_1_sva_10 <= cfg_lut_oflow_priority_1_sva_9;
      lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1 <= reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm
          & ({{22{lut_lookup_1_if_if_else_else_if_acc_itm_3}}, lut_lookup_1_if_if_else_else_if_acc_itm_3})
          & (signext_23_1(~ lut_lookup_1_if_if_else_acc_itm_9_1)) & (signext_23_1(~
          lut_lookup_if_if_lor_5_lpi_1_dfm_4));
      lut_lookup_le_fraction_1_lpi_1_dfm_22 <= (lut_lookup_if_else_else_else_else_mux_nl)
          & ({{34{lut_lookup_if_else_else_else_asn_mdf_1_sva_2}}, lut_lookup_if_else_else_else_asn_mdf_1_sva_2})
          & (signext_35_1(~ lut_lookup_if_else_else_slc_10_mdf_1_sva_4)) & ({{34{lut_lookup_1_if_else_slc_32_svs_8}},
          lut_lookup_1_if_else_slc_32_svs_8});
      lut_lookup_le_fraction_1_lpi_1_dfm_21 <= lut_lookup_1_else_else_else_else_rshift_itm
          & ({{34{lut_lookup_else_else_else_asn_mdf_1_sva_4}}, lut_lookup_else_else_else_asn_mdf_1_sva_4})
          & ({{34{lut_lookup_else_else_slc_32_mdf_1_sva_8}}, lut_lookup_else_else_slc_32_mdf_1_sva_8});
      lut_lookup_lo_fraction_1_lpi_1_dfm_9 <= lut_lookup_1_else_1_else_else_rshift_itm
          & (signext_35_1(~ lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3))
          & ({{34{lut_lookup_else_1_slc_32_mdf_1_sva_8}}, lut_lookup_else_1_slc_32_mdf_1_sva_8});
      lut_lookup_unequal_tmp_13 <= lut_lookup_else_unequal_tmp_18;
      lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1 <= reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg
          & ({{22{lut_lookup_2_if_if_else_else_if_acc_itm_3}}, lut_lookup_2_if_if_else_else_if_acc_itm_3})
          & (signext_23_1(~ lut_lookup_2_if_if_else_acc_itm_9_1)) & (signext_23_1(~
          lut_lookup_if_if_lor_6_lpi_1_dfm_4));
      lut_lookup_le_fraction_2_lpi_1_dfm_22 <= (lut_lookup_if_else_else_else_else_mux_1_nl)
          & ({{34{lut_lookup_if_else_else_else_asn_mdf_2_sva_2}}, lut_lookup_if_else_else_else_asn_mdf_2_sva_2})
          & (signext_35_1(~ lut_lookup_if_else_else_slc_10_mdf_2_sva_4)) & ({{34{lut_lookup_2_if_else_slc_32_svs_8}},
          lut_lookup_2_if_else_slc_32_svs_8});
      lut_lookup_le_fraction_2_lpi_1_dfm_21 <= lut_lookup_2_else_else_else_else_rshift_itm
          & ({{34{lut_lookup_else_else_else_asn_mdf_2_sva_4}}, lut_lookup_else_else_else_asn_mdf_2_sva_4})
          & ({{34{lut_lookup_else_else_slc_32_mdf_2_sva_8}}, lut_lookup_else_else_slc_32_mdf_2_sva_8});
      lut_lookup_lo_fraction_2_lpi_1_dfm_9 <= lut_lookup_2_else_1_else_else_rshift_itm
          & (signext_35_1(~ lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3))
          & ({{34{lut_lookup_else_1_slc_32_mdf_2_sva_8}}, lut_lookup_else_1_slc_32_mdf_2_sva_8});
      lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1 <= reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg
          & ({{22{lut_lookup_3_if_if_else_else_if_acc_itm_3}}, lut_lookup_3_if_if_else_else_if_acc_itm_3})
          & (signext_23_1(~ lut_lookup_3_if_if_else_acc_itm_9_1)) & (signext_23_1(~
          lut_lookup_if_if_lor_7_lpi_1_dfm_4));
      lut_lookup_le_fraction_3_lpi_1_dfm_22 <= (lut_lookup_if_else_else_else_else_mux_2_nl)
          & ({{34{lut_lookup_if_else_else_else_asn_mdf_3_sva_2}}, lut_lookup_if_else_else_else_asn_mdf_3_sva_2})
          & (signext_35_1(~ lut_lookup_if_else_else_slc_10_mdf_3_sva_4)) & ({{34{lut_lookup_3_if_else_slc_32_svs_8}},
          lut_lookup_3_if_else_slc_32_svs_8});
      lut_lookup_le_fraction_3_lpi_1_dfm_21 <= lut_lookup_3_else_else_else_else_rshift_itm
          & ({{34{lut_lookup_else_else_else_asn_mdf_3_sva_4}}, lut_lookup_else_else_else_asn_mdf_3_sva_4})
          & ({{34{lut_lookup_else_else_slc_32_mdf_3_sva_8}}, lut_lookup_else_else_slc_32_mdf_3_sva_8});
      lut_lookup_lo_fraction_3_lpi_1_dfm_9 <= lut_lookup_3_else_1_else_else_rshift_itm
          & (signext_35_1(~ lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3))
          & ({{34{lut_lookup_else_1_slc_32_mdf_3_sva_8}}, lut_lookup_else_1_slc_32_mdf_3_sva_8});
      lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1 <= reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1
          & ({{22{lut_lookup_4_if_if_else_else_if_acc_itm_3}}, lut_lookup_4_if_if_else_else_if_acc_itm_3})
          & (signext_23_1(~ lut_lookup_4_if_if_else_acc_itm_9_1)) & (signext_23_1(~
          lut_lookup_if_if_lor_1_lpi_1_dfm_4));
      lut_lookup_le_fraction_lpi_1_dfm_22 <= (lut_lookup_if_else_else_else_else_mux_3_nl)
          & ({{34{lut_lookup_if_else_else_else_asn_mdf_sva_2}}, lut_lookup_if_else_else_else_asn_mdf_sva_2})
          & (signext_35_1(~ lut_lookup_if_else_else_slc_10_mdf_sva_4)) & ({{34{lut_lookup_4_if_else_slc_32_svs_8}},
          lut_lookup_4_if_else_slc_32_svs_8});
      lut_lookup_le_fraction_lpi_1_dfm_21 <= lut_lookup_4_else_else_else_else_rshift_itm
          & ({{34{lut_lookup_else_else_else_asn_mdf_sva_4}}, lut_lookup_else_else_else_asn_mdf_sva_4})
          & ({{34{lut_lookup_else_else_slc_32_mdf_sva_8}}, lut_lookup_else_else_slc_32_mdf_sva_8});
      lut_lookup_lo_fraction_lpi_1_dfm_9 <= lut_lookup_4_else_1_else_else_rshift_itm
          & (signext_35_1(~ lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3))
          & ({{34{lut_lookup_else_1_slc_32_mdf_sva_8}}, lut_lookup_else_1_slc_32_mdf_sva_8});
      lut_in_data_sva_158 <= lut_in_data_sva_157;
      lut_lookup_1_and_svs_2 <= lut_lookup_else_mux_180_cse & lut_lookup_lo_uflow_1_lpi_1_dfm_3;
      lut_lookup_2_and_svs_2 <= lut_lookup_else_mux_182_cse & lut_lookup_lo_uflow_2_lpi_1_dfm_3;
      lut_lookup_3_and_svs_2 <= lut_lookup_else_mux_184_cse & lut_lookup_lo_uflow_3_lpi_1_dfm_3;
      cfg_lut_uflow_priority_1_sva_10 <= cfg_lut_uflow_priority_1_sva_9;
      lut_lookup_4_and_svs_2 <= lut_lookup_else_mux_186_cse & lut_lookup_lo_uflow_lpi_1_dfm_3;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_29 <= (lut_lookup_if_if_else_else_le_index_s_sva[5:0])
          & ({{5{lut_lookup_4_if_if_else_else_if_acc_itm_3}}, lut_lookup_4_if_if_else_else_if_acc_itm_3})
          & (signext_6_1(~ lut_lookup_4_if_if_else_acc_itm_9_1)) & (signext_6_1(~
          lut_lookup_if_if_lor_1_lpi_1_dfm_4));
      lut_lookup_le_index_0_5_0_lpi_1_dfm_28 <= lut_lookup_le_index_0_5_0_lpi_1_dfm_27;
      lut_lookup_le_index_0_5_0_lpi_1_dfm_26 <= lut_lookup_le_index_0_5_0_lpi_1_dfm_25;
      lut_lookup_else_unequal_tmp_13 <= lut_lookup_else_unequal_tmp_12;
      cfg_lut_le_function_1_sva_10 <= cfg_lut_le_function_1_sva_st_42;
      reg_lut_lookup_if_unequal_cse <= lut_lookup_if_unequal_tmp_1_mx0w0;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29 <= (lut_lookup_if_if_else_else_le_index_s_3_sva[5:0])
          & ({{5{lut_lookup_3_if_if_else_else_if_acc_itm_3}}, lut_lookup_3_if_if_else_else_if_acc_itm_3})
          & (signext_6_1(~ lut_lookup_3_if_if_else_acc_itm_9_1)) & (signext_6_1(~
          lut_lookup_if_if_lor_7_lpi_1_dfm_4));
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28 <= lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27;
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26 <= lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29 <= (lut_lookup_if_if_else_else_le_index_s_1_sva[5:0])
          & ({{5{lut_lookup_1_if_if_else_else_if_acc_itm_3}}, lut_lookup_1_if_if_else_else_if_acc_itm_3})
          & (signext_6_1(~ lut_lookup_1_if_if_else_acc_itm_9_1)) & (signext_6_1(~
          lut_lookup_if_if_lor_5_lpi_1_dfm_4));
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28 <= lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27;
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26 <= lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29 <= (lut_lookup_if_if_else_else_le_index_s_2_sva[5:0])
          & ({{5{lut_lookup_2_if_if_else_else_if_acc_itm_3}}, lut_lookup_2_if_if_else_else_if_acc_itm_3})
          & (signext_6_1(~ lut_lookup_2_if_if_else_acc_itm_9_1)) & (signext_6_1(~
          lut_lookup_if_if_lor_6_lpi_1_dfm_4));
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28 <= lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27;
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26 <= lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25;
      lut_lookup_lo_uflow_lpi_1_dfm_4 <= lut_lookup_lo_uflow_lpi_1_dfm_3;
      cfg_precision_1_sva_st_107 <= cfg_precision_1_sva_st_71;
      lut_lookup_lo_uflow_3_lpi_1_dfm_4 <= lut_lookup_lo_uflow_3_lpi_1_dfm_3;
      lut_lookup_lo_uflow_2_lpi_1_dfm_4 <= lut_lookup_lo_uflow_2_lpi_1_dfm_3;
      lut_lookup_lo_uflow_1_lpi_1_dfm_4 <= lut_lookup_lo_uflow_1_lpi_1_dfm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_2_else_else_if_mux_5_itm_1 <= 1'b0;
    end
    else if ( core_wen & (((mux_1139_nl) & or_cse) | lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1)
        ) begin
      lut_lookup_else_2_else_else_if_mux_5_itm_1 <= MUX_s_1_2_2(lut_lookup_lo_uflow_1_lpi_1_dfm_3,
          lut_lookup_else_mux_180_cse, lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_else_le_fra_1_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_267_nl) ) begin
      lut_lookup_else_if_else_le_fra_1_sva_4 <= lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_268_nl) ) begin
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_269_nl)) ) begin
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 <= IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_270_nl) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2 <= lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_5_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_274_nl)) ) begin
      lut_lookup_else_if_lor_5_lpi_1_dfm_6 <= lut_lookup_else_if_lor_5_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_5_lpi_1_dfm_st_3 <= 1'b0;
      lut_lookup_else_if_lor_7_lpi_1_dfm_st_3 <= 1'b0;
      lut_lookup_else_if_lor_1_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( lut_lookup_else_if_oelse_1_and_1_cse ) begin
      lut_lookup_else_if_lor_5_lpi_1_dfm_st_3 <= lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
      lut_lookup_else_if_lor_7_lpi_1_dfm_st_3 <= lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
      lut_lookup_else_if_lor_1_lpi_1_dfm_st_3 <= lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_72 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_276_nl) ) begin
      cfg_precision_1_sva_st_72 <= cfg_precision_1_sva_st_71;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_else_lo_fra_1_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_277_nl) ) begin
      lut_lookup_if_1_else_lo_fra_1_sva_4 <= lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_278_nl) ) begin
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_279_nl) ) begin
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 <= IsNaN_8U_23U_10_land_1_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_281_nl)) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2 <= lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_lor_5_lpi_1_dfm_5 <= 1'b0;
      lut_lookup_if_1_lor_6_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( lut_lookup_if_1_oelse_1_and_4_cse ) begin
      lut_lookup_if_1_lor_5_lpi_1_dfm_5 <= lut_lookup_if_1_lor_5_lpi_1_dfm_4;
      lut_lookup_if_1_lor_6_lpi_1_dfm_5 <= lut_lookup_if_1_lor_6_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_lor_5_lpi_1_dfm_st_4 <= 1'b0;
      lut_lookup_if_1_lor_6_lpi_1_dfm_st_4 <= 1'b0;
      lut_lookup_if_1_lor_7_lpi_1_dfm_st_4 <= 1'b0;
      lut_lookup_if_1_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( lut_lookup_if_1_oelse_1_and_5_cse ) begin
      lut_lookup_if_1_lor_5_lpi_1_dfm_st_4 <= lut_lookup_if_1_lor_5_lpi_1_dfm_4;
      lut_lookup_if_1_lor_6_lpi_1_dfm_st_4 <= lut_lookup_if_1_lor_6_lpi_1_dfm_4;
      lut_lookup_if_1_lor_7_lpi_1_dfm_st_4 <= lut_lookup_if_1_lor_7_lpi_1_dfm_4;
      lut_lookup_if_1_lor_1_lpi_1_dfm_st_4 <= lut_lookup_if_1_lor_1_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_2_else_else_if_mux_12_itm_1 <= 1'b0;
    end
    else if ( core_wen & (((mux_1152_nl) & or_cse) | lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1)
        ) begin
      lut_lookup_else_2_else_else_if_mux_12_itm_1 <= MUX_s_1_2_2(lut_lookup_lo_uflow_2_lpi_1_dfm_3,
          lut_lookup_else_mux_182_cse, lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_else_le_fra_2_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_286_nl) ) begin
      lut_lookup_else_if_else_le_fra_2_sva_4 <= lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_287_nl) ) begin
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_289_nl) ) begin
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 <= IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_291_nl) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2 <= lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_6_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_296_nl)) ) begin
      lut_lookup_else_if_lor_6_lpi_1_dfm_6 <= lut_lookup_else_if_lor_6_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_6_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_297_nl)) ) begin
      lut_lookup_else_if_lor_6_lpi_1_dfm_st_3 <= lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_else_lo_fra_2_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_299_nl) ) begin
      lut_lookup_if_1_else_lo_fra_2_sva_4 <= lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_300_nl) ) begin
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_301_nl)) ) begin
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 <= IsNaN_8U_23U_10_land_2_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_303_nl)) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2 <= lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_2_else_else_if_mux_19_itm_1 <= 1'b0;
    end
    else if ( core_wen & (((mux_1165_nl) & or_cse) | lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1)
        ) begin
      lut_lookup_else_2_else_else_if_mux_19_itm_1 <= MUX_s_1_2_2(lut_lookup_lo_uflow_3_lpi_1_dfm_3,
          lut_lookup_else_mux_184_cse, lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_else_le_fra_3_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_308_nl) ) begin
      lut_lookup_else_if_else_le_fra_3_sva_4 <= lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_309_nl) ) begin
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_310_nl)) ) begin
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 <= IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_311_nl) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2 <= lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_7_lpi_1_dfm_6 <= 1'b0;
      lut_lookup_else_if_lor_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( lut_lookup_else_if_oelse_1_and_4_cse ) begin
      lut_lookup_else_if_lor_7_lpi_1_dfm_6 <= lut_lookup_else_if_lor_7_lpi_1_dfm_5;
      lut_lookup_else_if_lor_1_lpi_1_dfm_6 <= lut_lookup_else_if_lor_1_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_else_lo_fra_3_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_319_nl) ) begin
      lut_lookup_if_1_else_lo_fra_3_sva_4 <= lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_320_nl)) ) begin
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_322_nl)) ) begin
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 <= IsNaN_8U_23U_10_land_3_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_325_nl)) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2 <= lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_lor_7_lpi_1_dfm_5 <= 1'b0;
      lut_lookup_if_1_lor_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( lut_lookup_if_1_oelse_1_and_8_cse ) begin
      lut_lookup_if_1_lor_7_lpi_1_dfm_5 <= lut_lookup_if_1_lor_7_lpi_1_dfm_4;
      lut_lookup_if_1_lor_1_lpi_1_dfm_5 <= lut_lookup_if_1_lor_1_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_2_else_else_if_mux_26_itm_1 <= 1'b0;
    end
    else if ( core_wen & (((mux_1178_nl) & or_cse) | lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1)
        ) begin
      lut_lookup_else_2_else_else_if_mux_26_itm_1 <= MUX_s_1_2_2(lut_lookup_lo_uflow_lpi_1_dfm_3,
          lut_lookup_else_mux_186_cse, lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_else_le_fra_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_332_nl) ) begin
      lut_lookup_else_if_else_le_fra_sva_4 <= lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_333_nl) ) begin
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2
          <= lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_334_nl)) ) begin
      IsNaN_8U_23U_6_land_lpi_1_dfm_7 <= IsNaN_8U_23U_6_land_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_335_nl) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2 <= lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_else_lo_fra_sva_4 <= 35'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_343_nl) ) begin
      lut_lookup_if_1_else_lo_fra_sva_4 <= lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_344_nl)) ) begin
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2
          <= lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_346_nl)) ) begin
      IsNaN_8U_23U_10_land_lpi_1_dfm_6 <= IsNaN_8U_23U_10_land_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2 <= 256'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_349_nl)) ) begin
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2 <= lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_le_uflow_lpi_1_dfm_6 <= 1'b0;
      lut_lookup_le_uflow_3_lpi_1_dfm_6 <= 1'b0;
      lut_lookup_le_uflow_2_lpi_1_dfm_6 <= 1'b0;
      lut_lookup_le_uflow_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( lut_lookup_le_uflow_and_cse ) begin
      lut_lookup_le_uflow_lpi_1_dfm_6 <= MUX_s_1_2_2(lut_lookup_else_mux_129_itm_2,
          lut_lookup_if_mux_123_mx0w1, and_dcpl_259);
      lut_lookup_le_uflow_3_lpi_1_dfm_6 <= MUX_s_1_2_2(lut_lookup_else_mux_86_itm_2,
          lut_lookup_if_mux_82_mx0w1, and_dcpl_259);
      lut_lookup_le_uflow_2_lpi_1_dfm_6 <= MUX_s_1_2_2(lut_lookup_else_mux_43_itm_2,
          lut_lookup_if_mux_41_mx0w1, and_dcpl_259);
      lut_lookup_le_uflow_1_lpi_1_dfm_6 <= MUX_s_1_2_2(lut_lookup_else_mux_itm_2,
          lut_lookup_if_mux_mx0w1, and_dcpl_259);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_13 <= 8'b0;
      lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2 <= 1'b0;
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13 <= 8'b0;
      lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2 <= 1'b0;
    end
    else if ( lut_lookup_lo_index_0_and_cse ) begin
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_13 <= lut_lookup_lo_index_0_7_0_lpi_1_dfm_12;
      lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2 <= lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          & lut_lookup_else_1_slc_32_mdf_sva_8;
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13 <= lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12;
      lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2 <= lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          & lut_lookup_else_1_slc_32_mdf_3_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 <= 1'b0;
      lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 <= 1'b0;
      lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 <= 1'b0;
    end
    else if ( lut_lookup_else_else_and_cse ) begin
      lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 <= MUX1HOT_s_1_3_2((lut_lookup_else_else_lut_lookup_else_else_and_10_nl),
          (lut_lookup_if_else_lut_lookup_if_else_and_11_nl), (lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_4_nl),
          {and_dcpl_258 , and_465_cse , and_466_cse});
      lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 <= MUX1HOT_s_1_3_2((lut_lookup_else_else_lut_lookup_else_else_and_7_nl),
          (lut_lookup_if_else_lut_lookup_if_else_and_12_nl), (lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_5_nl),
          {and_dcpl_258 , and_465_cse , and_466_cse});
      lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 <= MUX1HOT_s_1_3_2((lut_lookup_else_else_lut_lookup_else_else_and_4_nl),
          (lut_lookup_if_else_lut_lookup_if_else_and_13_nl), (lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_6_nl),
          {and_dcpl_258 , and_465_cse , and_466_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13 <= 8'b0;
      lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2 <= 1'b0;
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13 <= 8'b0;
      lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2 <= 1'b0;
    end
    else if ( lut_lookup_lo_index_0_and_2_cse ) begin
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13 <= lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12;
      lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2 <= lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          & lut_lookup_else_1_slc_32_mdf_2_sva_8;
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13 <= lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12;
      lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2 <= lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          & lut_lookup_else_1_slc_32_mdf_1_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_else_else_lut_lookup_else_else_or_3_cse & (mux_372_nl)
        ) begin
      lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 <= MUX1HOT_s_1_3_2((lut_lookup_else_else_lut_lookup_else_else_and_1_nl),
          (lut_lookup_if_else_lut_lookup_if_else_and_14_nl), (lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_7_nl),
          {and_dcpl_258 , and_465_cse , and_466_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_lo_uflow_1_lpi_1_dfm_3 <= 1'b0;
      lut_lookup_lo_uflow_2_lpi_1_dfm_3 <= 1'b0;
      lut_lookup_lo_uflow_3_lpi_1_dfm_3 <= 1'b0;
      lut_lookup_lo_uflow_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( lut_lookup_lo_uflow_and_4_cse ) begin
      lut_lookup_lo_uflow_1_lpi_1_dfm_3 <= MUX_s_1_2_2((~ lut_lookup_else_1_slc_32_mdf_1_sva_7),
          or_969_cse, and_636_cse);
      lut_lookup_lo_uflow_2_lpi_1_dfm_3 <= MUX_s_1_2_2((~ lut_lookup_else_1_slc_32_mdf_2_sva_7),
          lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0, and_636_cse);
      lut_lookup_lo_uflow_3_lpi_1_dfm_3 <= MUX_s_1_2_2((~ lut_lookup_else_1_slc_32_mdf_3_sva_7),
          lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0, and_636_cse);
      lut_lookup_lo_uflow_lpi_1_dfm_3 <= MUX_s_1_2_2((~ lut_lookup_else_1_slc_32_mdf_sva_7),
          lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0, and_636_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_1_and_46_cse ) begin
      FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[30:23]),
          (cfg_lut_le_start_rsci_d[30:23]), and_dcpl_280);
      FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3 <= readslicef_9_8_1((acc_4_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4 <= 8'b0;
      FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_2_and_44_cse ) begin
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[62:55]),
          (cfg_lut_lo_start_rsci_d[30:23]), and_dcpl_292);
      FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3 <= readslicef_9_8_1((acc_10_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4 <= 8'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_9_cse & (~ mux_tmp_4) ) begin
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[94:87]),
          (cfg_lut_lo_start_rsci_d[30:23]), and_dcpl_300);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_qr_lpi_1_dfm_4 <= 8'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_8_cse & (~ mux_tmp_4) ) begin
      FpAdd_8U_23U_2_qr_lpi_1_dfm_4 <= MUX_v_8_2_2((chn_lut_in_rsci_d_mxwt[126:119]),
          (cfg_lut_lo_start_rsci_d[30:23]), and_dcpl_308);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_a_greater_oelse_and_cse ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse,
          lut_lookup_1_else_else_acc_1_itm_32, and_dcpl_314);
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse,
          lut_lookup_2_else_else_acc_1_itm_32, and_dcpl_314);
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse,
          lut_lookup_3_else_else_acc_1_itm_32, and_dcpl_314);
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse,
          lut_lookup_4_else_else_acc_1_itm_32, and_dcpl_314);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_4_and_cse ) begin
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= MUX_s_1_2_2(lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1, and_dcpl_316);
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= MUX_s_1_2_2(lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1,
          lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0, and_dcpl_316);
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0, and_dcpl_315);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 <= 1'b0;
      FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 <= 1'b0;
      FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 <= 1'b0;
      FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_2_is_a_greater_oelse_and_cse ) begin
      FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse,
          lut_lookup_1_else_1_acc_itm_32, and_dcpl_314);
      FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse,
          lut_lookup_2_else_1_acc_itm_32, and_dcpl_314);
      FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse,
          lut_lookup_3_else_1_acc_itm_32, and_dcpl_314);
      FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse,
          lut_lookup_4_else_1_acc_itm_32, and_dcpl_314);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_4_and_1_cse ) begin
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= MUX_s_1_2_2(lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1, and_dcpl_316);
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= MUX_s_1_2_2(lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1,
          lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0, and_dcpl_316);
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= MUX_s_1_2_2(lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1, and_dcpl_316);
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= MUX_s_1_2_2(lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1,
          lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0, and_dcpl_316);
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= MUX_s_1_2_2(lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1, and_dcpl_316);
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= MUX_s_1_2_2(lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1,
          lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0, and_dcpl_316);
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0, and_dcpl_315);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ mux_582_itm) ) begin
      lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3 <= 8'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_9_cse & (~ mux_582_itm) ) begin
      FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3 <= readslicef_9_8_1((acc_9_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2 <= 1'b0;
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
    end
    else if ( IsZero_8U_23U_7_and_3_cse ) begin
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2 <= (cfg_lut_lo_start_rsci_d[30:0]!=31'b0000000000000000000000000000000);
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_a_right_shift_qr_sva_3 <= 8'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_8_cse & (~ mux_595_itm) ) begin
      FpAdd_8U_23U_2_a_right_shift_qr_sva_3 <= readslicef_9_8_1((acc_5_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_3_cse ) begin
      IsNaN_8U_23U_4_land_lpi_1_dfm_4 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2, and_524_rgt);
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_6,
          IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4, and_524_rgt);
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_6,
          IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4, and_524_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_4_cse ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_lpi_1_dfm_6,
          FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5, and_525_rgt);
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_1_land_1_lpi_1_dfm_6,
          FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5, and_525_rgt);
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4,
          FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4, and_525_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_5_cse ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_6,
          IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5,
          {and_527_rgt , and_529_rgt , and_525_rgt});
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_1_land_2_lpi_1_dfm_6,
          IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5,
          {and_527_rgt , and_529_rgt , and_525_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse & not_tmp_47
        ) begin
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 <= MUX_s_1_2_2(IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2, and_524_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_8U_23U_7_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_7_aelse_and_17_cse ) begin
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4,
          FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4, and_525_rgt);
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4,
          FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4, and_525_rgt);
      IsNaN_8U_23U_7_land_lpi_1_dfm_6 <= MUX_s_1_2_2(reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse,
          FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4, and_525_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_13_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_551_rgt | lut_lookup_or_17_rgt | lut_lookup_or_18_rgt)
        & not_tmp_47 ) begin
      FpAdd_8U_23U_1_mux_13_itm_3 <= MUX1HOT_s_1_3_2((lut_in_data_sva_154[31]), FpAdd_8U_23U_1_mux_1_itm_2,
          (~ (cfg_lut_le_start_1_sva_41[31])), {and_551_rgt , lut_lookup_or_17_rgt
          , lut_lookup_or_18_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_13_itm_1 <= 1'b0;
    end
    else if ( core_wen & (and_559_rgt | lut_lookup_and_126_rgt | lut_lookup_and_127_rgt
        | and_564_rgt) & (~ (mux_606_nl)) ) begin
      FpAdd_8U_23U_2_mux_13_itm_1 <= MUX1HOT_s_1_4_2((lut_in_data_sva_154[31]), FpAdd_8U_23U_2_mux_1_itm_2,
          (~ (cfg_lut_lo_start_1_sva_41[31])), FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0,
          {and_559_rgt , lut_lookup_and_126_rgt , lut_lookup_and_127_rgt , and_564_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_29_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_566_rgt | lut_lookup_and_124_rgt | lut_lookup_and_125_rgt)
        & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_1_mux_29_itm_3 <= MUX1HOT_s_1_3_2((lut_in_data_sva_154[63]), FpAdd_8U_23U_1_mux_17_itm_2,
          (~ (cfg_lut_le_start_1_sva_41[31])), {and_566_rgt , lut_lookup_and_124_rgt
          , lut_lookup_and_125_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_29_itm_1 <= 1'b0;
    end
    else if ( core_wen & (and_570_rgt | lut_lookup_and_122_rgt | lut_lookup_and_123_rgt
        | and_574_rgt) & (~ (mux_622_nl)) ) begin
      FpAdd_8U_23U_2_mux_29_itm_1 <= MUX1HOT_s_1_4_2((lut_in_data_sva_154[63]), FpAdd_8U_23U_2_mux_17_itm_2,
          (~ (cfg_lut_lo_start_1_sva_41[31])), FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0,
          {and_570_rgt , lut_lookup_and_122_rgt , lut_lookup_and_123_rgt , and_574_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_45_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_576_rgt | lut_lookup_and_120_rgt | lut_lookup_and_121_rgt)
        & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_1_mux_45_itm_3 <= MUX1HOT_s_1_3_2((lut_in_data_sva_154[95]), FpAdd_8U_23U_1_mux_33_itm_2,
          (~ (cfg_lut_le_start_1_sva_41[31])), {and_576_rgt , lut_lookup_and_120_rgt
          , lut_lookup_and_121_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_45_itm_1 <= 1'b0;
    end
    else if ( core_wen & (and_580_rgt | lut_lookup_and_118_rgt | lut_lookup_and_119_rgt
        | and_586_rgt) & (~ (mux_634_nl)) ) begin
      FpAdd_8U_23U_2_mux_45_itm_1 <= MUX1HOT_s_1_4_2((lut_in_data_sva_154[95]), FpAdd_8U_23U_2_mux_33_itm_2,
          (~ (cfg_lut_lo_start_1_sva_41[31])), FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0,
          {and_580_rgt , lut_lookup_and_118_rgt , lut_lookup_and_119_rgt , and_586_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_61_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_588_rgt | lut_lookup_or_rgt | lut_lookup_or_16_rgt)
        & (~ mux_25_itm) ) begin
      FpAdd_8U_23U_1_mux_61_itm_3 <= MUX1HOT_s_1_3_2((lut_in_data_sva_154[127]),
          FpAdd_8U_23U_1_mux_49_itm_2, (~ (cfg_lut_le_start_1_sva_41[31])), {and_588_rgt
          , lut_lookup_or_rgt , lut_lookup_or_16_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_61_itm_1 <= 1'b0;
    end
    else if ( core_wen & (and_595_rgt | lut_lookup_and_112_rgt | lut_lookup_and_113_rgt
        | and_586_rgt) & (~ (mux_651_nl)) ) begin
      FpAdd_8U_23U_2_mux_61_itm_1 <= MUX1HOT_s_1_4_2((lut_in_data_sva_154[127]),
          FpAdd_8U_23U_2_mux_49_itm_2, (~ (cfg_lut_lo_start_1_sva_41[31])), FpMantRNE_49U_24U_2_else_carry_sva_mx0w0,
          {and_595_rgt , lut_lookup_and_112_rgt , lut_lookup_and_113_rgt , and_586_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_1_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_653_nl) ) begin
      lut_lookup_else_else_else_le_index_u_1_sva_3 <= lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_1_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_654_nl) ) begin
      lut_lookup_else_1_lo_index_u_1_sva_3 <= nl_lut_lookup_else_1_lo_index_u_1_sva_3[31:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_2_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_655_nl) ) begin
      lut_lookup_else_else_else_le_index_u_2_sva_3 <= lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_2_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_657_nl) ) begin
      lut_lookup_else_1_lo_index_u_2_sva_3 <= nl_lut_lookup_else_1_lo_index_u_2_sva_3[31:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_3_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_658_nl) ) begin
      lut_lookup_else_else_else_le_index_u_3_sva_3 <= lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_3_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_659_nl) ) begin
      lut_lookup_else_1_lo_index_u_3_sva_3 <= nl_lut_lookup_else_1_lo_index_u_3_sva_3[31:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_660_nl) ) begin
      lut_lookup_else_else_else_le_index_u_sva_3 <= lut_lookup_if_else_else_le_data_sub_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_sva_3 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_661_nl) ) begin
      lut_lookup_else_1_lo_index_u_sva_3 <= nl_lut_lookup_else_1_lo_index_u_sva_3[31:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse & (mux_667_nl)
        ) begin
      IsNaN_8U_23U_6_land_lpi_1_dfm_6 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp,
          lut_lookup_4_if_else_else_else_else_acc_itm_32_1, FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6,
          lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3, {and_604_rgt , and_606_rgt , and_dcpl_403
          , and_dcpl_405});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_1_lpi_1_dfm_5 <= 1'b0;
      lut_lookup_else_if_lor_7_lpi_1_dfm_5 <= 1'b0;
      lut_lookup_else_if_lor_6_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( lut_lookup_else_if_oelse_1_and_8_cse ) begin
      lut_lookup_else_if_lor_1_lpi_1_dfm_5 <= lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1;
      lut_lookup_else_if_lor_7_lpi_1_dfm_5 <= lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1;
      lut_lookup_else_if_lor_6_lpi_1_dfm_5 <= lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_unequal_tmp_12 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_672_nl) ) begin
      lut_lookup_else_unequal_tmp_12 <= lut_lookup_unequal_tmp_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse & (mux_678_nl)
        ) begin
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp,
          lut_lookup_3_if_else_else_else_else_acc_itm_32_1, FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6,
          lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3, {and_604_rgt , and_606_rgt , and_dcpl_403
          , and_dcpl_405});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse & (mux_689_nl)
        ) begin
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp,
          lut_lookup_2_if_else_else_else_else_acc_itm_32_1, FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6,
          lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3, {and_604_rgt , and_606_rgt , and_dcpl_403
          , and_dcpl_405});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse & (mux_700_nl)
        ) begin
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 <= MUX1HOT_s_1_4_2(and_1142_cse, lut_lookup_1_if_else_else_else_else_acc_itm_32_1,
          FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6, lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3,
          {and_604_rgt , and_606_rgt , and_dcpl_403 , and_dcpl_405});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_if_lor_5_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_704_nl)) ) begin
      lut_lookup_else_if_lor_5_lpi_1_dfm_5 <= lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_12 <= 8'b0;
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12 <= 8'b0;
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= 1'b0;
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= 1'b0;
    end
    else if ( lut_lookup_lo_index_0_and_4_cse ) begin
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_12 <= lut_lookup_lo_index_0_7_0_lpi_1_dfm_11;
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12 <= lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11;
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse & (mux_711_nl)
        ) begin
      IsNaN_8U_23U_10_land_lpi_1_dfm_5 <= MUX_s_1_2_2(and_1138_cse, FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5,
          and_427_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_lor_1_lpi_1_dfm_4 <= 1'b0;
      lut_lookup_if_1_lor_7_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( lut_lookup_if_1_oelse_1_and_12_cse ) begin
      lut_lookup_if_1_lor_1_lpi_1_dfm_4 <= lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0;
      lut_lookup_if_1_lor_7_lpi_1_dfm_4 <= lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse & (mux_722_nl)
        ) begin
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 <= MUX_s_1_2_2(and_1139_cse, FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5,
          and_427_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12 <= 8'b0;
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12 <= 8'b0;
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= 1'b0;
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= 1'b0;
    end
    else if ( lut_lookup_lo_index_0_and_6_cse ) begin
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12 <= lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11;
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12 <= lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11;
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4
          <= lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse & (mux_732_nl)
        ) begin
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 <= MUX_s_1_2_2(and_1140_cse, FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5,
          and_427_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_1_lor_6_lpi_1_dfm_4 <= 1'b0;
      lut_lookup_if_1_lor_5_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( lut_lookup_if_1_oelse_1_and_14_cse ) begin
      lut_lookup_if_1_lor_6_lpi_1_dfm_4 <= lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0;
      lut_lookup_if_1_lor_5_lpi_1_dfm_4 <= or_969_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse & (mux_739_nl)
        ) begin
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 <= MUX_s_1_2_2(and_1141_cse, FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5,
          and_427_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_if_lor_5_lpi_1_dfm_4 <= 1'b0;
      lut_lookup_if_if_lor_6_lpi_1_dfm_4 <= 1'b0;
      lut_lookup_if_if_lor_7_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( lut_lookup_if_if_oelse_1_and_cse ) begin
      lut_lookup_if_if_lor_5_lpi_1_dfm_4 <= lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3;
      lut_lookup_if_if_lor_6_lpi_1_dfm_4 <= lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3;
      lut_lookup_if_if_lor_7_lpi_1_dfm_4 <= lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_else_asn_mdf_1_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_759_nl) ) begin
      lut_lookup_if_else_else_else_asn_mdf_1_sva_2 <= lut_lookup_1_if_else_else_else_if_acc_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_1_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_768_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_1_sva_4 <= lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_if_else_slc_32_svs_8 <= 1'b0;
      lut_lookup_2_if_else_slc_32_svs_8 <= 1'b0;
      lut_lookup_3_if_else_slc_32_svs_8 <= 1'b0;
    end
    else if ( lut_lookup_if_else_if_and_4_cse ) begin
      lut_lookup_1_if_else_slc_32_svs_8 <= lut_lookup_1_if_else_slc_32_svs_7;
      lut_lookup_2_if_else_slc_32_svs_8 <= lut_lookup_2_if_else_slc_32_svs_7;
      lut_lookup_3_if_else_slc_32_svs_8 <= lut_lookup_3_if_else_slc_32_svs_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm <= 8'b0;
    end
    else if ( and_dcpl_648 & (~ cfg_lut_le_function_1_sva_st_41) & or_1857_cse &
        lut_lookup_1_if_else_slc_32_svs_7 & (~ lut_lookup_if_else_else_slc_10_mdf_1_sva_3)
        & FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & lut_lookup_1_if_else_else_else_if_acc_itm_3
        & (~(nor_874_cse | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8)) ) begin
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm <= IntLog2_32U_mux1h_1_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm <= 23'b0;
    end
    else if ( (mux_1246_nl) & and_dcpl_648 & or_cse ) begin
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm <= IntLog2_32U_mux1h_1_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_783_nl) ) begin
      lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[1:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_8 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_784_nl) ) begin
      cfg_precision_1_sva_8 <= cfg_precision_1_sva_st_70;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_else_else_else_else_le_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_785_nl) ) begin
      lut_lookup_1_else_else_else_else_le_data_f_and_itm_2 <= lut_lookup_else_else_else_le_index_u_1_sva_4
          & lut_lookup_1_else_else_else_else_le_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_else_else_else_else_acc_reg <= 1'b0;
      reg_lut_lookup_2_else_else_else_else_acc_reg <= 1'b0;
      reg_lut_lookup_3_else_else_else_else_acc_reg <= 1'b0;
      reg_lut_lookup_4_else_else_else_else_acc_reg <= 1'b0;
    end
    else if ( and_898_cse ) begin
      reg_lut_lookup_1_else_else_else_else_acc_reg <= lut_lookup_else_else_else_else_mux1h_rgt[8];
      reg_lut_lookup_2_else_else_else_else_acc_reg <= lut_lookup_else_else_else_else_mux1h_1_rgt[8];
      reg_lut_lookup_3_else_else_else_else_acc_reg <= lut_lookup_else_else_else_else_mux1h_2_rgt[8];
      reg_lut_lookup_4_else_else_else_else_acc_reg <= lut_lookup_else_else_else_else_mux1h_3_rgt[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_else_else_else_else_acc_1_reg <= 1'b0;
      reg_lut_lookup_2_else_else_else_else_acc_1_reg <= 1'b0;
      reg_lut_lookup_3_else_else_else_else_acc_1_reg <= 1'b0;
      reg_lut_lookup_4_else_else_else_else_acc_1_reg <= 1'b0;
    end
    else if ( and_901_cse ) begin
      reg_lut_lookup_1_else_else_else_else_acc_1_reg <= lut_lookup_else_else_else_else_mux1h_rgt[7];
      reg_lut_lookup_2_else_else_else_else_acc_1_reg <= lut_lookup_else_else_else_else_mux1h_1_rgt[7];
      reg_lut_lookup_3_else_else_else_else_acc_1_reg <= lut_lookup_else_else_else_else_mux1h_2_rgt[7];
      reg_lut_lookup_4_else_else_else_else_acc_1_reg <= lut_lookup_else_else_else_else_mux1h_3_rgt[7];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_else_else_else_else_acc_2_reg <= 3'b0;
    end
    else if ( (and_896_cse | cfg_lut_le_function_1_sva_st_41 | (~ lut_lookup_1_if_else_else_else_else_acc_itm_32_1))
        & or_cse & core_wen ) begin
      reg_lut_lookup_1_else_else_else_else_acc_2_reg <= lut_lookup_else_else_else_else_mux1h_rgt[6:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_else_else_else_else_acc_3_reg <= 4'b0;
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg <= 23'b0;
      reg_lut_lookup_2_else_else_else_else_acc_3_reg <= 4'b0;
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg <= 23'b0;
      reg_lut_lookup_3_else_else_else_else_acc_3_reg <= 4'b0;
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 <= 23'b0;
      reg_lut_lookup_4_else_else_else_else_acc_3_reg <= 4'b0;
    end
    else if ( and_905_cse ) begin
      reg_lut_lookup_1_else_else_else_else_acc_3_reg <= lut_lookup_else_else_else_else_mux1h_rgt[3:0];
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg <= IntLog2_32U_IntLog2_32U_mux_rgt[22:0];
      reg_lut_lookup_2_else_else_else_else_acc_3_reg <= lut_lookup_else_else_else_else_mux1h_1_rgt[3:0];
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg <= IntLog2_32U_IntLog2_32U_mux_1_rgt[22:0];
      reg_lut_lookup_3_else_else_else_else_acc_3_reg <= lut_lookup_else_else_else_else_mux1h_2_rgt[3:0];
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 <= IntLog2_32U_IntLog2_32U_mux_2_rgt[22:0];
      reg_lut_lookup_4_else_else_else_else_acc_3_reg <= lut_lookup_else_else_else_else_mux1h_3_rgt[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_1_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_792_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_1_sva_4 <= lut_lookup_else_else_else_asn_mdf_1_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_slc_32_mdf_1_sva_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_797_nl) ) begin
      lut_lookup_else_else_slc_32_mdf_1_sva_8 <= lut_lookup_else_else_slc_32_mdf_1_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 <= 23'b0;
    end
    else if ( core_wen & ((or_cse & IsNaN_8U_23U_7_land_1_lpi_1_dfm_7) | and_653_rgt)
        & (~ (mux_798_nl)) ) begin
      FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 <= MUX_v_23_2_2((lut_in_data_sva_156[22:0]),
          FpAdd_8U_23U_2_asn_50_mx0w1, and_653_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_799_nl)) ) begin
      lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2 <= lut_lookup_else_1_lo_index_u_1_sva_4
          & lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_else_1_else_else_acc_itm <= 1'b0;
    end
    else if ( core_wen & (~ FpAdd_8U_23U_2_mux_13_itm_3) & main_stage_v_3 & or_1857_cse
        & lut_lookup_else_1_slc_32_mdf_1_sva_7 & (~ FpMantRNE_49U_24U_2_else_carry_1_sva_2)
        & FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 & or_cse ) begin
      reg_lut_lookup_1_else_1_else_else_acc_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_1_else_1_else_else_acc_1_itm <= 8'b0;
    end
    else if ( (~ (mux_1248_nl)) & core_wen & (~ FpAdd_8U_23U_2_mux_13_itm_3) & main_stage_v_3
        & or_cse ) begin
      reg_lut_lookup_1_else_1_else_else_acc_1_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_803_nl) ) begin
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= FpMantRNE_49U_24U_2_else_carry_1_sva_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_806_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_8 <= lut_lookup_else_1_slc_32_mdf_1_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_else_asn_mdf_2_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_823_nl) ) begin
      lut_lookup_if_else_else_else_asn_mdf_2_sva_2 <= lut_lookup_2_if_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_2_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_832_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_2_sva_4 <= lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg <= 8'b0;
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg <= 8'b0;
      reg_IntLog2_32U_ac_int_cctor_1_30_0_reg <= 8'b0;
    end
    else if ( and_907_cse ) begin
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg <= IntLog2_32U_IntLog2_32U_mux_rgt[30:23];
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg <= IntLog2_32U_IntLog2_32U_mux_1_rgt[30:23];
      reg_IntLog2_32U_ac_int_cctor_1_30_0_reg <= IntLog2_32U_IntLog2_32U_mux_2_rgt[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_840_nl) ) begin
      lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[1:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_else_else_else_else_le_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_841_nl) ) begin
      lut_lookup_2_else_else_else_else_le_data_f_and_itm_2 <= lut_lookup_else_else_else_le_index_u_2_sva_4
          & lut_lookup_1_else_else_else_else_le_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_2_else_else_else_else_acc_2_reg <= 3'b0;
    end
    else if ( (and_896_cse | cfg_lut_le_function_1_sva_st_41 | (~ lut_lookup_2_if_else_else_else_else_acc_itm_32_1))
        & or_cse & core_wen ) begin
      reg_lut_lookup_2_else_else_else_else_acc_2_reg <= lut_lookup_else_else_else_else_mux1h_1_rgt[6:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_2_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_848_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_2_sva_4 <= lut_lookup_else_else_else_asn_mdf_2_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_slc_32_mdf_2_sva_8 <= 1'b0;
      lut_lookup_else_else_slc_32_mdf_3_sva_8 <= 1'b0;
      lut_lookup_else_else_slc_32_mdf_sva_8 <= 1'b0;
    end
    else if ( lut_lookup_else_else_and_5_cse ) begin
      lut_lookup_else_else_slc_32_mdf_2_sva_8 <= lut_lookup_else_else_slc_32_mdf_2_sva_7;
      lut_lookup_else_else_slc_32_mdf_3_sva_8 <= lut_lookup_else_else_slc_32_mdf_3_sva_7;
      lut_lookup_else_else_slc_32_mdf_sva_8 <= lut_lookup_else_else_slc_32_mdf_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 <= 23'b0;
    end
    else if ( core_wen & ((or_cse & IsNaN_8U_23U_7_land_2_lpi_1_dfm_7) | and_661_rgt)
        & (~ (mux_854_nl)) ) begin
      FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 <= MUX_v_23_2_2((lut_in_data_sva_156[54:32]),
          FpAdd_8U_23U_2_asn_45_mx0w1, and_661_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_855_nl)) ) begin
      lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2 <= lut_lookup_else_1_lo_index_u_2_sva_4
          & lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_2_else_1_else_else_acc_itm <= 1'b0;
    end
    else if ( core_wen & (~ FpAdd_8U_23U_2_mux_29_itm_3) & main_stage_v_3 & or_1857_cse
        & lut_lookup_else_1_slc_32_mdf_2_sva_7 & (~ FpMantRNE_49U_24U_2_else_carry_2_sva_2)
        & FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 & or_cse ) begin
      reg_lut_lookup_2_else_1_else_else_acc_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_2_else_1_else_else_acc_1_itm <= 8'b0;
    end
    else if ( (~ (mux_1250_nl)) & core_wen & (~ FpAdd_8U_23U_2_mux_29_itm_3) & main_stage_v_3
        & or_cse ) begin
      reg_lut_lookup_2_else_1_else_else_acc_1_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_859_nl) ) begin
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= FpMantRNE_49U_24U_2_else_carry_2_sva_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_2_sva_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_861_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_2_sva_8 <= lut_lookup_else_1_slc_32_mdf_2_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_else_asn_mdf_3_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_878_nl) ) begin
      lut_lookup_if_else_else_else_asn_mdf_3_sva_2 <= lut_lookup_3_if_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_3_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_887_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_3_sva_4 <= lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_895_nl) ) begin
      lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[1:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_else_else_else_else_le_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_896_nl) ) begin
      lut_lookup_3_else_else_else_else_le_data_f_and_itm_2 <= lut_lookup_else_else_else_le_index_u_3_sva_4
          & lut_lookup_1_else_else_else_else_le_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_3_else_else_else_else_acc_2_reg <= 3'b0;
    end
    else if ( (and_896_cse | cfg_lut_le_function_1_sva_st_41 | (~ lut_lookup_3_if_else_else_else_else_acc_itm_32_1))
        & or_cse & core_wen ) begin
      reg_lut_lookup_3_else_else_else_else_acc_2_reg <= lut_lookup_else_else_else_else_mux1h_2_rgt[6:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_3_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_903_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_3_sva_4 <= lut_lookup_else_else_else_asn_mdf_3_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 <= 23'b0;
    end
    else if ( core_wen & ((or_cse & IsNaN_8U_23U_7_land_3_lpi_1_dfm_7) | and_668_rgt)
        & (~ (mux_910_nl)) ) begin
      FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 <= MUX_v_23_2_2((lut_in_data_sva_156[86:64]),
          FpAdd_8U_23U_2_asn_40_mx0w1, and_668_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_912_nl)) ) begin
      lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2 <= lut_lookup_else_1_lo_index_u_3_sva_4
          & lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_3_else_1_else_else_acc_itm <= 1'b0;
    end
    else if ( core_wen & (~ FpAdd_8U_23U_2_mux_45_itm_3) & main_stage_v_3 & or_1857_cse
        & lut_lookup_else_1_slc_32_mdf_3_sva_7 & (~ FpMantRNE_49U_24U_2_else_carry_3_sva_2)
        & FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 & or_cse ) begin
      reg_lut_lookup_3_else_1_else_else_acc_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_3_else_1_else_else_acc_1_itm <= 8'b0;
    end
    else if ( (mux_1251_nl) & core_wen & (~ FpAdd_8U_23U_2_mux_45_itm_3) & main_stage_v_3
        & or_cse ) begin
      reg_lut_lookup_3_else_1_else_else_acc_1_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_916_nl) ) begin
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= FpMantRNE_49U_24U_2_else_carry_3_sva_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_3_sva_8 <= 1'b0;
      lut_lookup_else_1_slc_32_mdf_sva_8 <= 1'b0;
    end
    else if ( lut_lookup_else_1_and_6_cse ) begin
      lut_lookup_else_1_slc_32_mdf_3_sva_8 <= lut_lookup_else_1_slc_32_mdf_3_sva_7;
      lut_lookup_else_1_slc_32_mdf_sva_8 <= lut_lookup_else_1_slc_32_mdf_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_if_lor_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_926_nl) ) begin
      lut_lookup_if_if_lor_1_lpi_1_dfm_4 <= lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_else_asn_mdf_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_936_nl) ) begin
      lut_lookup_if_else_else_else_asn_mdf_sva_2 <= lut_lookup_4_if_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_slc_10_mdf_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_945_nl) ) begin
      lut_lookup_if_else_else_slc_10_mdf_sva_4 <= lut_lookup_if_else_else_slc_10_mdf_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_if_else_slc_32_svs_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_953_nl) ) begin
      lut_lookup_4_if_else_slc_32_svs_8 <= lut_lookup_4_if_else_slc_32_svs_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_954_nl) ) begin
      lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3
          <= reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[1:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_else_else_else_else_le_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_955_nl) ) begin
      lut_lookup_4_else_else_else_else_le_data_f_and_itm_2 <= lut_lookup_else_else_else_le_index_u_sva_4
          & lut_lookup_1_else_else_else_else_le_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_4_else_else_else_else_acc_2_reg <= 3'b0;
    end
    else if ( (and_896_cse | cfg_lut_le_function_1_sva_st_41 | (~ lut_lookup_4_if_else_else_else_else_acc_itm_32_1))
        & or_cse & core_wen ) begin
      reg_lut_lookup_4_else_else_else_else_acc_2_reg <= lut_lookup_else_else_else_else_mux1h_3_rgt[6:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_962_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_sva_4 <= lut_lookup_else_else_else_asn_mdf_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 <= 23'b0;
    end
    else if ( core_wen & ((or_cse & IsNaN_8U_23U_7_land_lpi_1_dfm_7) | and_676_rgt)
        & (~ (mux_969_nl)) ) begin
      FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 <= MUX_v_23_2_2((lut_in_data_sva_156[118:96]),
          FpAdd_8U_23U_2_asn_35_mx0w1, and_676_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_971_nl)) ) begin
      lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2 <= lut_lookup_else_1_lo_index_u_sva_4
          & lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_4_else_1_else_else_acc_itm <= 1'b0;
    end
    else if ( core_wen & (~ FpAdd_8U_23U_2_mux_61_itm_3) & main_stage_v_3 & or_1857_cse
        & lut_lookup_else_1_slc_32_mdf_sva_7 & (~ FpMantRNE_49U_24U_2_else_carry_sva_2)
        & FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 & or_cse ) begin
      reg_lut_lookup_4_else_1_else_else_acc_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_lut_lookup_4_else_1_else_else_acc_1_itm <= 8'b0;
    end
    else if ( (mux_1252_nl) & core_wen & (~ FpAdd_8U_23U_2_mux_61_itm_3) & main_stage_v_3
        & or_cse ) begin
      reg_lut_lookup_4_else_1_else_else_acc_1_itm <= lut_lookup_else_1_else_else_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_975_nl) ) begin
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
          <= FpMantRNE_49U_24U_2_else_carry_sva_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_mux_129_itm_2 <= 1'b0;
      lut_lookup_else_mux_86_itm_2 <= 1'b0;
      lut_lookup_else_mux_43_itm_2 <= 1'b0;
    end
    else if ( lut_lookup_else_and_8_cse ) begin
      lut_lookup_else_mux_129_itm_2 <= MUX_s_1_2_2((~ lut_lookup_else_else_slc_32_mdf_sva_7),
          lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1, and_636_cse);
      lut_lookup_else_mux_86_itm_2 <= MUX_s_1_2_2((~ lut_lookup_else_else_slc_32_mdf_3_sva_7),
          lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1, and_636_cse);
      lut_lookup_else_mux_43_itm_2 <= MUX_s_1_2_2((~ lut_lookup_else_else_slc_32_mdf_2_sva_7),
          lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1, and_636_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_mux_itm_2 <= 1'b0;
    end
    else if ( core_wen & (and_427_cse | and_679_rgt) & mux_tmp_978 ) begin
      lut_lookup_else_mux_itm_2 <= MUX_s_1_2_2((~ lut_lookup_else_else_slc_32_mdf_1_sva_7),
          lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1, and_679_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_981_nl) ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2 <= lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_slc_32_mdf_1_sva_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_986_nl) ) begin
      lut_lookup_else_else_slc_32_mdf_1_sva_7 <= lut_lookup_1_if_else_slc_32_svs_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_1_sva_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_995_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_1_sva_3 <= lut_lookup_1_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_997_nl) ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1 <= lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_slc_32_mdf_2_sva_7 <= 1'b0;
      lut_lookup_else_else_slc_32_mdf_3_sva_7 <= 1'b0;
      lut_lookup_else_else_slc_32_mdf_sva_7 <= 1'b0;
    end
    else if ( lut_lookup_else_else_and_9_cse ) begin
      lut_lookup_else_else_slc_32_mdf_2_sva_7 <= lut_lookup_2_if_else_slc_32_svs_6;
      lut_lookup_else_else_slc_32_mdf_3_sva_7 <= lut_lookup_3_if_else_slc_32_svs_6;
      lut_lookup_else_else_slc_32_mdf_sva_7 <= lut_lookup_4_if_else_slc_32_svs_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_2_sva_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1013_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_2_sva_3 <= lut_lookup_2_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1015_nl) ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1 <= lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_3_sva_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1031_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_3_sva_3 <= lut_lookup_3_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_sva_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1033_nl) ) begin
      IntLog2_32U_ac_int_cctor_1_30_0_sva_1 <= lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_asn_mdf_sva_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1049_nl) ) begin
      lut_lookup_else_else_else_asn_mdf_sva_3 <= lut_lookup_4_else_else_else_if_acc_itm_3_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_sva_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1051_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_sva_7 <= lut_lookup_else_1_slc_32_mdf_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_3_sva_7 <= 1'b0;
      lut_lookup_else_1_slc_32_mdf_2_sva_7 <= 1'b0;
    end
    else if ( lut_lookup_else_1_and_9_cse ) begin
      lut_lookup_else_1_slc_32_mdf_3_sva_7 <= lut_lookup_else_1_slc_32_mdf_3_sva_6;
      lut_lookup_else_1_slc_32_mdf_2_sva_7 <= lut_lookup_else_1_slc_32_mdf_2_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1055_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_7 <= lut_lookup_else_1_slc_32_mdf_1_sva_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_11 <= 8'b0;
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11 <= 8'b0;
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11 <= 8'b0;
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11 <= 8'b0;
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= 1'b0;
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= 1'b0;
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= 1'b0;
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= 1'b0;
    end
    else if ( lut_lookup_lo_index_0_and_8_cse ) begin
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_11 <= (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0])
          & (signext_8_1(~ (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])))
          & ({{7{lut_lookup_else_1_slc_32_mdf_sva_6}}, lut_lookup_else_1_slc_32_mdf_sva_6});
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11 <= (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0])
          & (signext_8_1(~ (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])))
          & ({{7{lut_lookup_else_1_slc_32_mdf_3_sva_6}}, lut_lookup_else_1_slc_32_mdf_3_sva_6});
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11 <= (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0])
          & (signext_8_1(~ (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])))
          & ({{7{lut_lookup_else_1_slc_32_mdf_2_sva_6}}, lut_lookup_else_1_slc_32_mdf_2_sva_6});
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11 <= (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0])
          & (signext_8_1(~ (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])))
          & ({{7{lut_lookup_else_1_slc_32_mdf_1_sva_6}}, lut_lookup_else_1_slc_32_mdf_1_sva_6});
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3
          <= lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_1_or_11_cse & (mux_1058_nl) ) begin
      FpAdd_8U_23U_1_mux_1_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[31]), (~
          (cfg_lut_le_start_rsci_d[31])), and_dcpl_280);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_nor_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1059_nl) ) begin
      IsNaN_8U_23U_4_nor_itm_2 <= IsNaN_8U_23U_4_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2 <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse & (mux_1060_nl)
        ) begin
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2 <= MUX_s_1_2_2(IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0,
          IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0, and_dcpl_316);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1061_nl) ) begin
      FpAdd_8U_23U_2_mux_1_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[31]), (~
          (cfg_lut_lo_start_rsci_d[31])), and_dcpl_284);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_17_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1062_nl) ) begin
      FpAdd_8U_23U_1_mux_17_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[63]), (~
          (cfg_lut_le_start_rsci_d[31])), and_dcpl_288);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_17_itm_2 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_10_cse & (mux_1063_nl) ) begin
      FpAdd_8U_23U_2_mux_17_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[63]), (~
          (cfg_lut_lo_start_rsci_d[31])), and_dcpl_292);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_33_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1064_nl) ) begin
      FpAdd_8U_23U_1_mux_33_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[95]), (~
          (cfg_lut_le_start_rsci_d[31])), and_dcpl_296);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_33_itm_2 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_9_cse & (mux_1066_nl) ) begin
      FpAdd_8U_23U_2_mux_33_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[95]), (~
          (cfg_lut_lo_start_rsci_d[31])), and_dcpl_300);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_8_nor_2_itm_2 <= 1'b0;
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_8_and_cse ) begin
      IsNaN_8U_23U_8_nor_2_itm_2 <= IsNaN_8U_23U_8_nor_2_tmp_1;
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2 <= IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_mux_49_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1069_nl) ) begin
      FpAdd_8U_23U_1_mux_49_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[127]), (~
          (cfg_lut_le_start_rsci_d[31])), and_dcpl_304);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_nor_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1070_nl) ) begin
      IsNaN_8U_23U_4_nor_3_itm_2 <= IsNaN_8U_23U_4_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse & (mux_1071_nl)
        ) begin
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2 <= MUX_s_1_2_2(IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0,
          IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0, and_dcpl_316);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_2_mux_49_itm_2 <= 1'b0;
    end
    else if ( core_wen & lut_lookup_FpAdd_8U_23U_2_or_8_cse & (mux_1073_nl) ) begin
      FpAdd_8U_23U_2_mux_49_itm_2 <= MUX_s_1_2_2((chn_lut_in_rsci_d_mxwt[127]), (~
          (cfg_lut_lo_start_rsci_d[31])), and_dcpl_308);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_8_nor_3_itm_2 <= 1'b0;
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_8_and_2_cse ) begin
      IsNaN_8U_23U_8_nor_3_itm_2 <= IsNaN_8U_23U_8_nor_2_tmp_1;
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2 <= IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= 6'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse & (mux_1077_nl)
        ) begin
      lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= MUX_v_6_2_2((lut_lookup_if_else_else_else_le_index_s_1_sva[5:0]), (lut_lookup_else_else_else_lut_lookup_else_else_else_and_1_nl),
          and_dcpl_148);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_1_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1078_nl) ) begin
      lut_lookup_else_else_else_le_index_u_1_sva_4 <= lut_lookup_else_else_else_le_index_u_1_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_1_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_1079_nl)) ) begin
      lut_lookup_else_1_lo_index_u_1_sva_4 <= lut_lookup_else_1_lo_index_u_1_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= 6'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse & (mux_1084_nl)
        ) begin
      lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= MUX_v_6_2_2((lut_lookup_if_else_else_else_le_index_s_2_sva[5:0]), (lut_lookup_else_else_else_lut_lookup_else_else_else_and_3_nl),
          and_dcpl_148);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_2_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1085_nl) ) begin
      lut_lookup_else_else_else_le_index_u_2_sva_4 <= lut_lookup_else_else_else_le_index_u_2_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_2_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_1086_nl)) ) begin
      lut_lookup_else_1_lo_index_u_2_sva_4 <= lut_lookup_else_1_lo_index_u_2_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= 6'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse & (mux_1091_nl)
        ) begin
      lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= MUX_v_6_2_2((lut_lookup_if_else_else_else_le_index_s_3_sva[5:0]), (lut_lookup_else_else_else_lut_lookup_else_else_else_and_5_nl),
          and_dcpl_148);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_3_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1092_nl) ) begin
      lut_lookup_else_else_else_le_index_u_3_sva_4 <= lut_lookup_else_else_else_le_index_u_3_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_3_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_1093_nl)) ) begin
      lut_lookup_else_1_lo_index_u_3_sva_4 <= lut_lookup_else_1_lo_index_u_3_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= 6'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse & (mux_1096_nl)
        ) begin
      lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2
          <= MUX_v_6_2_2((lut_lookup_if_else_else_else_le_index_s_sva[5:0]), (lut_lookup_else_else_else_lut_lookup_else_else_else_and_7_nl),
          and_dcpl_148);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_else_else_le_index_u_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1097_nl) ) begin
      lut_lookup_else_else_else_le_index_u_sva_4 <= lut_lookup_else_else_else_le_index_u_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_lo_index_u_sva_4 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_1098_nl)) ) begin
      lut_lookup_else_1_lo_index_u_sva_4 <= lut_lookup_else_1_lo_index_u_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (~ (mux_1101_nl)) ) begin
      lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1 <= lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1103_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_6 <= lut_lookup_else_1_slc_32_mdf_1_sva_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1104_nl) ) begin
      lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1 <= lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_2_sva_6 <= 1'b0;
      lut_lookup_else_1_slc_32_mdf_3_sva_6 <= 1'b0;
    end
    else if ( lut_lookup_else_1_and_13_cse ) begin
      lut_lookup_else_1_slc_32_mdf_2_sva_6 <= lut_lookup_else_1_slc_32_mdf_2_sva_5;
      lut_lookup_else_1_slc_32_mdf_3_sva_6 <= lut_lookup_else_1_slc_32_mdf_3_sva_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1107_nl) ) begin
      lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1 <= lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1110_nl) ) begin
      lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1 <= lut_lookup_if_else_else_le_data_sub_sva_mx0w0[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_sva_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1112_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_sva_6 <= lut_lookup_else_1_slc_32_mdf_sva_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_sva_5 <= 1'b0;
      lut_lookup_else_1_slc_32_mdf_3_sva_5 <= 1'b0;
      lut_lookup_else_1_slc_32_mdf_2_sva_5 <= 1'b0;
    end
    else if ( lut_lookup_else_1_and_16_cse ) begin
      lut_lookup_else_1_slc_32_mdf_sva_5 <= lut_lookup_4_else_1_acc_itm_32;
      lut_lookup_else_1_slc_32_mdf_3_sva_5 <= lut_lookup_3_else_1_acc_itm_32;
      lut_lookup_else_1_slc_32_mdf_2_sva_5 <= lut_lookup_2_else_1_acc_itm_32;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_5 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_54) & (mux_1118_nl) ) begin
      lut_lookup_else_1_slc_32_mdf_1_sva_5 <= lut_lookup_1_else_1_acc_itm_32;
    end
  end
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_7_nl = MUX1HOT_v_12_5_2((lut_lookup_le_fraction_1_lpi_1_dfm_22[11:0]),
      (lut_lookup_le_fraction_1_lpi_1_dfm_9[11:0]), (lut_lookup_le_fraction_1_lpi_1_dfm_21[11:0]),
      (lut_lookup_lo_fraction_1_lpi_1_dfm_1[11:0]), (lut_lookup_lo_fraction_1_lpi_1_dfm_9[11:0]),
      {lut_lookup_and_5_cse , lut_lookup_and_6_cse , lut_lookup_and_7_cse , lut_lookup_and_138_cse
      , lut_lookup_and_139_cse});
  assign lut_lookup_not_39_nl = ~ lut_lookup_lut_lookup_nor_19_cse;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_6_nl = MUX1HOT_v_12_5_2((lut_lookup_le_fraction_2_lpi_1_dfm_22[11:0]),
      (lut_lookup_le_fraction_2_lpi_1_dfm_9[11:0]), (lut_lookup_le_fraction_2_lpi_1_dfm_21[11:0]),
      (lut_lookup_lo_fraction_2_lpi_1_dfm_1[11:0]), (lut_lookup_lo_fraction_2_lpi_1_dfm_9[11:0]),
      {lut_lookup_and_13_cse , lut_lookup_and_14_cse , lut_lookup_and_15_cse , lut_lookup_and_136_cse
      , lut_lookup_and_137_cse});
  assign lut_lookup_not_38_nl = ~ lut_lookup_lut_lookup_nor_18_cse;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_5_nl = MUX1HOT_v_12_5_2((lut_lookup_le_fraction_3_lpi_1_dfm_22[11:0]),
      (lut_lookup_le_fraction_3_lpi_1_dfm_9[11:0]), (lut_lookup_le_fraction_3_lpi_1_dfm_21[11:0]),
      (lut_lookup_lo_fraction_3_lpi_1_dfm_1[11:0]), (lut_lookup_lo_fraction_3_lpi_1_dfm_9[11:0]),
      {lut_lookup_and_21_cse , lut_lookup_and_22_cse , lut_lookup_and_23_cse , lut_lookup_and_134_cse
      , lut_lookup_and_135_cse});
  assign lut_lookup_not_37_nl = ~ lut_lookup_lut_lookup_nor_17_cse;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_4_nl = MUX1HOT_v_12_5_2((lut_lookup_le_fraction_lpi_1_dfm_22[11:0]),
      (lut_lookup_le_fraction_lpi_1_dfm_9[11:0]), (lut_lookup_le_fraction_lpi_1_dfm_21[11:0]),
      (lut_lookup_lo_fraction_lpi_1_dfm_1[11:0]), (lut_lookup_lo_fraction_lpi_1_dfm_9[11:0]),
      {lut_lookup_and_29_cse , lut_lookup_and_30_cse , lut_lookup_and_31_cse , lut_lookup_and_132_cse
      , lut_lookup_and_133_cse});
  assign lut_lookup_not_36_nl = ~ lut_lookup_lut_lookup_nor_16_cse;
  assign lut_lookup_else_2_if_mux_5_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0, cfg_lut_oflow_priority_1_sva_10);
  assign lut_lookup_else_2_else_else_mux_61_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0, cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_nl = (lut_lookup_else_2_else_else_mux_61_nl)
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse;
  assign lut_lookup_else_2_mux_1_nl = MUX_s_1_2_2((lut_lookup_else_2_else_lut_lookup_else_2_else_and_nl),
      (lut_lookup_else_2_if_mux_5_nl), lut_lookup_1_else_2_and_svs);
  assign lut_lookup_else_2_if_mux_11_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0, cfg_lut_oflow_priority_1_sva_10);
  assign lut_lookup_else_2_else_else_mux_60_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0, cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_2_nl = (lut_lookup_else_2_else_else_mux_60_nl)
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse;
  assign lut_lookup_else_2_mux_27_nl = MUX_s_1_2_2((lut_lookup_else_2_else_lut_lookup_else_2_else_and_2_nl),
      (lut_lookup_else_2_if_mux_11_nl), lut_lookup_2_else_2_and_svs);
  assign lut_lookup_else_2_if_mux_17_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0, cfg_lut_oflow_priority_1_sva_10);
  assign lut_lookup_else_2_else_else_mux_59_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0, cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_4_nl = (lut_lookup_else_2_else_else_mux_59_nl)
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse;
  assign lut_lookup_else_2_mux_53_nl = MUX_s_1_2_2((lut_lookup_else_2_else_lut_lookup_else_2_else_and_4_nl),
      (lut_lookup_else_2_if_mux_17_nl), lut_lookup_3_else_2_and_svs);
  assign lut_lookup_else_2_if_mux_23_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0, cfg_lut_oflow_priority_1_sva_10);
  assign lut_lookup_else_2_else_else_mux_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0,
      lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0, cfg_lut_hybrid_priority_1_sva_10);
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_6_nl = (lut_lookup_else_2_else_else_mux_nl)
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse;
  assign lut_lookup_else_2_mux_79_nl = MUX_s_1_2_2((lut_lookup_else_2_else_lut_lookup_else_2_else_and_6_nl),
      (lut_lookup_else_2_if_mux_23_nl), lut_lookup_4_else_2_and_svs);
  assign lut_lookup_else_if_lut_lookup_else_if_and_2_nl = (lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1[5:0])
      & ({{5{lut_lookup_1_else_if_else_if_acc_itm_3_1}}, lut_lookup_1_else_if_else_if_acc_itm_3_1})
      & (signext_6_1(~ lut_lookup_else_if_lor_5_lpi_1_dfm_6));
  assign lut_lookup_else_if_lut_lookup_else_if_and_5_nl = (lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1[5:0])
      & ({{5{lut_lookup_2_else_if_else_if_acc_itm_3_1}}, lut_lookup_2_else_if_else_if_acc_itm_3_1})
      & (signext_6_1(~ lut_lookup_else_if_lor_6_lpi_1_dfm_6));
  assign lut_lookup_else_if_lut_lookup_else_if_and_8_nl = (lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1[5:0])
      & ({{5{lut_lookup_3_else_if_else_if_acc_itm_3_1}}, lut_lookup_3_else_if_else_if_acc_itm_3_1})
      & (signext_6_1(~ lut_lookup_else_if_lor_7_lpi_1_dfm_6));
  assign lut_lookup_else_if_lut_lookup_else_if_and_11_nl = (lut_lookup_else_if_else_le_int_lpi_1_dfm_1[5:0])
      & ({{5{lut_lookup_4_else_if_else_if_acc_itm_3_1}}, lut_lookup_4_else_if_else_if_acc_itm_3_1})
      & (signext_6_1(~ lut_lookup_else_if_lor_1_lpi_1_dfm_6));
  assign lut_lookup_else_2_lut_lookup_else_2_and_4_nl = lut_lookup_else_2_else_else_if_mux_5_itm_1
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse
      & (~ lut_lookup_1_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_3_nl = MUX_s_1_2_2(lut_lookup_le_miss_1_sva,
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse);
  assign lut_lookup_else_2_else_mux_3_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_3_nl),
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_103_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_3_nl),
      cfg_lut_oflow_priority_1_sva_10, lut_lookup_1_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_13_nl = MUX_s_1_2_2(z_out, lut_lookup_else_2_else_if_mux_2_cse_mx0,
      lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse);
  assign lut_lookup_else_2_else_mux_18_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_13_nl),
      lut_lookup_else_2_else_if_mux_2_cse_mx0, lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_107_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_18_nl),
      z_out, lut_lookup_1_else_2_and_svs);
  assign lut_lookup_if_2_mux_21_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_uflow_priority_1_sva_10);
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_1_nl = (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_3_nl
      = (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1]) & lut_lookup_le_miss_1_sva;
  assign lut_lookup_else_2_else_else_mux_12_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_3_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse);
  assign lut_lookup_else_2_else_mux_17_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_12_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse, lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_108_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_17_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_1_nl), lut_lookup_1_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_8_nl = (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_nl = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_2_nl
      = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 & lut_lookup_le_miss_1_sva;
  assign lut_lookup_else_2_else_else_mux_11_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_2_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse);
  assign lut_lookup_else_2_else_mux_16_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_11_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse, lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_109_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_16_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_nl), lut_lookup_1_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_9_nl = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_lut_lookup_else_2_and_5_nl = lut_lookup_else_2_else_else_if_mux_12_itm_1
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse
      & (~ lut_lookup_2_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_18_nl = MUX_s_1_2_2(lut_lookup_le_miss_2_sva,
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse);
  assign lut_lookup_else_2_else_mux_23_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_18_nl),
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_104_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_23_nl),
      cfg_lut_oflow_priority_1_sva_10, lut_lookup_2_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_28_nl = MUX_s_1_2_2(z_out_1, lut_lookup_else_2_else_if_mux_7_cse_mx0,
      lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse);
  assign lut_lookup_else_2_else_mux_38_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_28_nl),
      lut_lookup_else_2_else_if_mux_7_cse_mx0, lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_110_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_38_nl),
      z_out_1, lut_lookup_2_else_2_and_svs);
  assign lut_lookup_if_2_mux_22_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_uflow_priority_1_sva_10);
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_3_nl = (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_7_nl
      = (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1]) & lut_lookup_le_miss_2_sva;
  assign lut_lookup_else_2_else_else_mux_27_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_7_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse);
  assign lut_lookup_else_2_else_mux_37_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_27_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse, lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_111_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_37_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_3_nl), lut_lookup_2_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_10_nl = (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_2_nl = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_6_nl
      = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 & lut_lookup_le_miss_2_sva;
  assign lut_lookup_else_2_else_else_mux_26_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_6_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse);
  assign lut_lookup_else_2_else_mux_36_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_26_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse, lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_112_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_36_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_2_nl), lut_lookup_2_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_11_nl = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_lut_lookup_else_2_and_6_nl = lut_lookup_else_2_else_else_if_mux_19_itm_1
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse
      & (~ lut_lookup_3_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_33_nl = MUX_s_1_2_2(lut_lookup_le_miss_3_sva,
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse);
  assign lut_lookup_else_2_else_mux_43_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_33_nl),
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_105_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_43_nl),
      cfg_lut_oflow_priority_1_sva_10, lut_lookup_3_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_43_nl = MUX_s_1_2_2(z_out_2, lut_lookup_else_2_else_if_mux_12_cse_mx0,
      lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse);
  assign lut_lookup_else_2_else_mux_58_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_43_nl),
      lut_lookup_else_2_else_if_mux_12_cse_mx0, lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_113_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_58_nl),
      z_out_2, lut_lookup_3_else_2_and_svs);
  assign lut_lookup_if_2_mux_23_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_uflow_priority_1_sva_10);
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_5_nl = (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_11_nl
      = (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1]) & lut_lookup_le_miss_3_sva;
  assign lut_lookup_else_2_else_else_mux_42_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_11_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse);
  assign lut_lookup_else_2_else_mux_57_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_42_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse, lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_114_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_57_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_5_nl), lut_lookup_3_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_12_nl = (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_4_nl = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_10_nl
      = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 & lut_lookup_le_miss_3_sva;
  assign lut_lookup_else_2_else_else_mux_41_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_10_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse);
  assign lut_lookup_else_2_else_mux_56_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_41_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse, lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_115_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_56_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_4_nl), lut_lookup_3_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_13_nl = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_lut_lookup_else_2_and_7_nl = lut_lookup_else_2_else_else_if_mux_26_itm_1
      & lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse
      & (~ lut_lookup_4_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_48_nl = MUX_s_1_2_2(lut_lookup_le_miss_sva,
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse);
  assign lut_lookup_else_2_else_mux_63_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_48_nl),
      cfg_lut_hybrid_priority_1_sva_10, lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_106_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_63_nl),
      cfg_lut_oflow_priority_1_sva_10, lut_lookup_4_else_2_and_svs);
  assign lut_lookup_else_2_else_else_mux_58_nl = MUX_s_1_2_2(z_out_3, lut_lookup_else_2_else_if_mux_17_cse_mx0,
      lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse);
  assign lut_lookup_else_2_else_mux_78_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_58_nl),
      lut_lookup_else_2_else_if_mux_17_cse_mx0, lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_116_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_78_nl),
      z_out_3, lut_lookup_4_else_2_and_svs);
  assign lut_lookup_if_2_mux_24_nl = MUX_s_1_2_2(lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0,
      (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[0]), cfg_lut_uflow_priority_1_sva_10);
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_7_nl = (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_15_nl
      = (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1]) & lut_lookup_le_miss_sva;
  assign lut_lookup_else_2_else_else_mux_57_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_15_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse);
  assign lut_lookup_else_2_else_mux_77_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_57_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse, lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_117_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_77_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_7_nl), lut_lookup_4_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_14_nl = (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1])
      & cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_6_nl = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0
      & cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_14_nl
      = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 & lut_lookup_le_miss_sva;
  assign lut_lookup_else_2_else_else_mux_56_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_14_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse, lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse);
  assign lut_lookup_else_2_else_mux_76_nl = MUX_s_1_2_2((lut_lookup_else_2_else_else_mux_56_nl),
      lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse, lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs);
  assign lut_lookup_else_2_mux_118_nl = MUX_s_1_2_2((lut_lookup_else_2_else_mux_76_nl),
      (lut_lookup_else_2_if_lut_lookup_else_2_if_and_6_nl), lut_lookup_4_else_2_and_svs);
  assign lut_lookup_if_2_lut_lookup_if_2_and_15_nl = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0
      & cfg_lut_uflow_priority_1_sva_10;
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_10_nl = MUX_v_8_2_2((cfg_lut_lo_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[30:23]), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1);
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_11_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[30:23])),
      (~ (cfg_lut_lo_start_rsci_d[30:23])), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1);
  assign nl_acc_6_nl = ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_10_nl) , 1'b1})
      + ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_11_nl) , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[8:0];
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_12_nl = MUX_v_8_2_2((cfg_lut_le_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[62:55]), FpAdd_8U_23U_b_right_shift_qif_and_tmp_2);
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_13_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[62:55])),
      (~ (cfg_lut_le_start_rsci_d[30:23])), FpAdd_8U_23U_b_right_shift_qif_and_tmp_2);
  assign nl_acc_8_nl = ({(FpAdd_8U_23U_a_right_shift_qelse_mux_12_nl) , 1'b1}) +
      ({(FpAdd_8U_23U_a_right_shift_qelse_mux_13_nl) , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[8:0];
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_14_nl = MUX_v_8_2_2((cfg_lut_le_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[94:87]), FpAdd_8U_23U_b_right_shift_qif_and_tmp_3);
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_15_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[94:87])),
      (~ (cfg_lut_le_start_rsci_d[30:23])), FpAdd_8U_23U_b_right_shift_qif_and_tmp_3);
  assign nl_acc_11_nl = ({(FpAdd_8U_23U_a_right_shift_qelse_mux_14_nl) , 1'b1}) +
      ({(FpAdd_8U_23U_a_right_shift_qelse_mux_15_nl) , 1'b1});
  assign acc_11_nl = nl_acc_11_nl[8:0];
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_10_nl = MUX_v_8_2_2((cfg_lut_le_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[126:119]), FpAdd_8U_23U_b_right_shift_qif_and_tmp_1);
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_11_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[126:119])),
      (~ (cfg_lut_le_start_rsci_d[30:23])), FpAdd_8U_23U_b_right_shift_qif_and_tmp_1);
  assign nl_acc_7_nl = ({(FpAdd_8U_23U_a_right_shift_qelse_mux_10_nl) , 1'b1}) +
      ({(FpAdd_8U_23U_a_right_shift_qelse_mux_11_nl) , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[8:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl[49:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl[49:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl[49:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl[49:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl[49:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl[49:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl[49:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl[49:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl[49:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl[49:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl[49:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl[49:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0);
  assign lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl[49:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0);
  assign lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl[49:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0);
  assign lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl[49:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0) + 50'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl[49:0];
  assign mux_1209_nl = MUX_s_1_2_2(or_1689_cse, (~ main_stage_v_2), IsNaN_8U_23U_1_land_1_lpi_1_dfm_7);
  assign mux_13_nl = MUX_s_1_2_2((mux_1209_nl), or_1689_cse, reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign mux_1210_nl = MUX_s_1_2_2(or_tmp_63, (~ main_stage_v_3), FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6);
  assign mux_38_nl = MUX_s_1_2_2((mux_1210_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign mux_39_nl = MUX_s_1_2_2((mux_38_nl), (mux_13_nl), or_cse);
  assign or_2081_nl = nor_874_cse | or_tmp_1663;
  assign or_1931_nl = (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_1_sva_3
      | (~ lut_lookup_1_if_else_slc_32_svs_7);
  assign mux_1218_nl = MUX_s_1_2_2((or_1931_nl), or_tmp_1663, or_cse);
  assign nor_793_nl = ~(nor_792_cse | cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6));
  assign mux_1219_nl = MUX_s_1_2_2((mux_1218_nl), (or_2081_nl), nor_793_nl);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl = MUX_v_2_2_2(2'b00, (lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt[7:6]),
      FpNormalize_8U_49U_oelse_not_9);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl = MUX_v_6_2_2(6'b000000,
      (lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt[5:0]), FpNormalize_8U_49U_oelse_not_9);
  assign mux_1125_nl = MUX_s_1_2_2(and_896_cse, or_dcpl_51, or_cse);
  assign FpAdd_8U_23U_o_expo_or_3_nl = FpAdd_8U_23U_and_51_ssc | (~ (mux_1125_nl));
  assign or_1941_nl = (reg_cfg_precision_1_sva_st_13_cse_1[0]) | (~((reg_cfg_precision_1_sva_st_13_cse_1[1])
      & or_1936_cse));
  assign mux_1222_nl = MUX_s_1_2_2(or_tmp_1671, (~ or_1936_cse), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_1223_nl = MUX_s_1_2_2((mux_1222_nl), or_tmp_1671, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign mux_1224_nl = MUX_s_1_2_2((mux_1223_nl), (or_1941_nl), lut_lookup_1_if_else_else_acc_itm_10);
  assign and_868_nl = reg_cfg_lut_le_function_1_sva_st_20_cse & IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign mux_57_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, and_868_nl);
  assign and_869_nl = cfg_lut_le_function_1_sva_st_41 & FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign mux_58_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, and_869_nl);
  assign mux_59_nl = MUX_s_1_2_2((mux_58_nl), (mux_57_nl), or_cse);
  assign nor_772_nl = ~(IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 | or_tmp_101);
  assign nor_773_nl = ~(IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 | FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5
      | IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 | (~
      main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign mux_61_nl = MUX_s_1_2_2((nor_773_nl), (nor_772_nl), or_cse);
  assign nor_769_nl = ~(IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 | nor_13_cse | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5
      | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 | (~ main_stage_v_2));
  assign mux_62_nl = MUX_s_1_2_2(nor_tmp_12, (nor_769_nl), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_63_nl = MUX_s_1_2_2((mux_62_nl), nor_tmp_12, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign nor_770_nl = ~(IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 | FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5);
  assign mux_64_nl = MUX_s_1_2_2(nor_tmp_14, (nor_770_nl), cfg_precision_1_sva_st_70[1]);
  assign mux_65_nl = MUX_s_1_2_2((mux_64_nl), nor_tmp_14, cfg_precision_1_sva_st_70[0]);
  assign and_45_nl = main_stage_v_3 & (mux_65_nl);
  assign mux_66_nl = MUX_s_1_2_2((and_45_nl), (mux_63_nl), or_cse);
  assign nl_lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl = FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)})
      + 8'b1;
  assign lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl = nl_lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_nl = MUX_v_8_2_2(8'b00000000,
      (lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl), FpNormalize_8U_49U_2_oelse_not_9);
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5
      + 8'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl = nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0];
  assign or_114_nl = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6
      | or_tmp_101;
  assign mux_67_nl = MUX_s_1_2_2((or_114_nl), or_1689_cse, lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp);
  assign or_118_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 | (~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10);
  assign mux_68_nl = MUX_s_1_2_2((or_118_nl), or_tmp_63, lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign mux_69_nl = MUX_s_1_2_2((mux_68_nl), (mux_67_nl), or_cse);
  assign mux_74_nl = MUX_s_1_2_2(mux_tmp_72, (~ main_stage_v_2), IsNaN_8U_23U_8_land_lpi_1_dfm_4);
  assign or_120_nl = (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10) | IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  assign mux_75_nl = MUX_s_1_2_2((mux_74_nl), mux_tmp_72, or_120_nl);
  assign mux_80_nl = MUX_s_1_2_2(mux_tmp_78, (~ main_stage_v_3), IsNaN_8U_23U_8_land_2_lpi_1_dfm_7);
  assign or_125_nl = (cfg_precision_1_sva_st_70!=2'b10) | IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign mux_81_nl = MUX_s_1_2_2((mux_80_nl), mux_tmp_78, or_125_nl);
  assign mux_82_nl = MUX_s_1_2_2((mux_81_nl), (mux_75_nl), or_cse);
  assign mux_84_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, IsNaN_8U_23U_7_land_1_lpi_1_dfm_6);
  assign mux_85_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5);
  assign mux_86_nl = MUX_s_1_2_2((mux_85_nl), (mux_84_nl), or_cse);
  assign or_40_nl = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) | reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_23_nl = MUX_s_1_2_2((~ main_stage_v_2), or_1689_cse, or_40_nl);
  assign mux_87_nl = MUX_s_1_2_2(or_tmp_63, (~ main_stage_v_3), FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6);
  assign mux_88_nl = MUX_s_1_2_2((mux_87_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign mux_89_nl = MUX_s_1_2_2((mux_88_nl), (mux_23_nl), or_cse);
  assign or_2080_nl = nor_874_cse | or_tmp_1674;
  assign or_1948_nl = (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_2_sva_3
      | (~ lut_lookup_2_if_else_slc_32_svs_7);
  assign mux_1225_nl = MUX_s_1_2_2((or_1948_nl), or_tmp_1674, or_cse);
  assign nor_796_nl = ~(nor_792_cse | cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6));
  assign mux_1226_nl = MUX_s_1_2_2((mux_1225_nl), (or_2080_nl), nor_796_nl);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl = MUX_v_2_2_2(2'b00, (lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt[7:6]),
      FpNormalize_8U_49U_oelse_not_11);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_10_nl = MUX_v_6_2_2(6'b000000,
      (lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt[5:0]), FpNormalize_8U_49U_oelse_not_11);
  assign FpAdd_8U_23U_o_expo_or_2_nl = FpAdd_8U_23U_and_53_ssc | (~ mux_1126_cse);
  assign nor_852_nl = ~(lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp | nor_855_cse);
  assign mux_1229_nl = MUX_s_1_2_2(or_tmp_1678, (nor_852_nl), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_1230_nl = MUX_s_1_2_2((mux_1229_nl), or_tmp_1678, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign and_864_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_119_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, and_864_nl);
  assign and_865_nl = cfg_lut_le_function_1_sva_st_41 & FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign mux_120_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, and_865_nl);
  assign mux_121_nl = MUX_s_1_2_2((mux_120_nl), (mux_119_nl), or_cse);
  assign nor_760_nl = ~(nor_31_cse | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10)
      | IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 | IsNaN_8U_23U_7_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6);
  assign nor_761_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10) |
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6
      | FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5);
  assign mux_123_nl = MUX_s_1_2_2((nor_761_nl), (nor_760_nl), or_cse);
  assign nor_757_nl = ~(IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 | nor_31_cse | IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5
      | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 | (~ main_stage_v_2));
  assign mux_124_nl = MUX_s_1_2_2(nor_tmp_32, (nor_757_nl), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_125_nl = MUX_s_1_2_2((mux_124_nl), nor_tmp_32, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign nor_758_nl = ~(IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6 | FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5);
  assign mux_126_nl = MUX_s_1_2_2(nor_tmp_34, (nor_758_nl), cfg_precision_1_sva_st_70[1]);
  assign mux_127_nl = MUX_s_1_2_2((mux_126_nl), nor_tmp_34, cfg_precision_1_sva_st_70[0]);
  assign and_48_nl = main_stage_v_3 & (mux_127_nl);
  assign mux_128_nl = MUX_s_1_2_2((and_48_nl), (mux_125_nl), or_cse);
  assign nl_lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl = FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)})
      + 8'b1;
  assign lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl = nl_lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_2_nl = MUX_v_8_2_2(8'b00000000,
      (lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl), FpNormalize_8U_49U_2_oelse_not_11);
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5
      + 8'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl = nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0];
  assign and_49_nl = or_cse & mux_tmp_128;
  assign or_184_nl = (~(IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_7
      | FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5)) | lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign mux_130_nl = MUX_s_1_2_2(nand_tmp_4, (and_49_nl), or_184_nl);
  assign nor_35_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10));
  assign mux_131_nl = MUX_s_1_2_2(nand_tmp_4, (mux_130_nl), nor_35_nl);
  assign mux_133_nl = MUX_s_1_2_2((~ or_tmp_44), main_stage_v_2, IsNaN_8U_23U_7_land_2_lpi_1_dfm_6);
  assign mux_134_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5);
  assign mux_135_nl = MUX_s_1_2_2((mux_134_nl), (mux_133_nl), or_cse);
  assign mux_27_nl = MUX_s_1_2_2((~ main_stage_v_2), or_1689_cse, or_48_cse);
  assign mux_1211_nl = MUX_s_1_2_2(or_tmp_63, (~ main_stage_v_3), FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6);
  assign mux_137_nl = MUX_s_1_2_2((mux_1211_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign mux_138_nl = MUX_s_1_2_2((mux_137_nl), (mux_27_nl), or_cse);
  assign or_2079_nl = nor_874_cse | or_tmp_1684;
  assign or_1964_nl = (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_3_sva_3
      | (~ lut_lookup_3_if_else_slc_32_svs_7);
  assign mux_1231_nl = MUX_s_1_2_2((or_1964_nl), or_tmp_1684, or_cse);
  assign nor_799_nl = ~(nor_792_cse | cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6));
  assign mux_1232_nl = MUX_s_1_2_2((mux_1231_nl), (or_2079_nl), nor_799_nl);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl = MUX_v_2_2_2(2'b00, (lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt[7:6]),
      FpNormalize_8U_49U_oelse_not_13);
  assign mux_1233_nl = MUX_s_1_2_2(IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5, IsNaN_8U_23U_4_land_3_lpi_1_dfm_5,
      reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl = MUX_v_6_2_2(6'b000000,
      (lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt[5:0]), FpNormalize_8U_49U_oelse_not_13);
  assign FpAdd_8U_23U_o_expo_or_1_nl = FpAdd_8U_23U_and_55_ssc | (~ mux_1126_cse);
  assign or_1976_nl = (reg_cfg_precision_1_sva_st_13_cse_1[0]) | (~((reg_cfg_precision_1_sva_st_13_cse_1[1])
      & or_tmp_1692));
  assign mux_1235_nl = MUX_s_1_2_2(or_48_cse, (~ or_tmp_1692), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_1236_nl = MUX_s_1_2_2((mux_1235_nl), or_48_cse, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign mux_1237_nl = MUX_s_1_2_2((mux_1236_nl), (or_1976_nl), lut_lookup_3_if_else_else_acc_itm_10);
  assign and_861_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_155_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, and_861_nl);
  assign and_862_nl = cfg_lut_le_function_1_sva_st_41 & FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign mux_156_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, and_862_nl);
  assign mux_157_nl = MUX_s_1_2_2((mux_156_nl), (mux_155_nl), or_cse);
  assign nor_745_nl = ~(IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 | nor_42_cse | IsNaN_8U_23U_7_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10));
  assign nor_746_nl = ~(IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 | FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5
      | IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 | IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 | (cfg_precision_1_sva_st_70!=2'b10)
      | (~ main_stage_v_3));
  assign mux_159_nl = MUX_s_1_2_2((nor_746_nl), (nor_745_nl), or_cse);
  assign nor_742_nl = ~(IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 | nor_42_cse | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5
      | IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 | (~ main_stage_v_2));
  assign mux_160_nl = MUX_s_1_2_2(nor_tmp_44, (nor_742_nl), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_161_nl = MUX_s_1_2_2((mux_160_nl), nor_tmp_44, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign nor_743_nl = ~(IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_3_lpi_1_dfm_5
      | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 | FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5);
  assign mux_162_nl = MUX_s_1_2_2(nor_tmp_46, (nor_743_nl), cfg_precision_1_sva_st_70[1]);
  assign mux_163_nl = MUX_s_1_2_2((mux_162_nl), nor_tmp_46, cfg_precision_1_sva_st_70[0]);
  assign and_54_nl = main_stage_v_3 & (mux_163_nl);
  assign mux_164_nl = MUX_s_1_2_2((and_54_nl), (mux_161_nl), or_cse);
  assign nl_lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl = FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17)})
      + 8'b1;
  assign lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl = nl_lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_4_nl = MUX_v_8_2_2(8'b00000000,
      (lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl), FpNormalize_8U_49U_2_oelse_not_13);
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5
      + 8'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl = nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0];
  assign or_247_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 | nor_42_cse | IsNaN_8U_23U_7_land_3_lpi_1_dfm_6
      | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10);
  assign mux_165_nl = MUX_s_1_2_2((or_247_nl), or_1689_cse, lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp);
  assign or_251_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 | IsNaN_8U_23U_8_land_3_lpi_1_dfm_5
      | IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 | (cfg_precision_1_sva_st_70!=2'b10) |
      (~ main_stage_v_3);
  assign mux_166_nl = MUX_s_1_2_2((or_251_nl), or_tmp_63, lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2);
  assign mux_167_nl = MUX_s_1_2_2((mux_166_nl), (mux_165_nl), or_cse);
  assign mux_169_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, IsNaN_8U_23U_7_land_3_lpi_1_dfm_6);
  assign mux_170_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5);
  assign mux_171_nl = MUX_s_1_2_2((mux_170_nl), (mux_169_nl), or_cse);
  assign mux_31_nl = MUX_s_1_2_2(or_1689_cse, (~ main_stage_v_2), IsNaN_8U_23U_1_land_lpi_1_dfm_7);
  assign mux_32_nl = MUX_s_1_2_2((mux_31_nl), or_1689_cse, reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign mux_1212_nl = MUX_s_1_2_2(or_tmp_63, (~ main_stage_v_3), FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6);
  assign mux_173_nl = MUX_s_1_2_2((mux_1212_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign mux_174_nl = MUX_s_1_2_2((mux_173_nl), (mux_32_nl), or_cse);
  assign or_2078_nl = nor_874_cse | or_tmp_1697;
  assign or_1983_nl = (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_sva_3
      | (~ lut_lookup_4_if_else_slc_32_svs_7);
  assign mux_1238_nl = MUX_s_1_2_2((or_1983_nl), or_tmp_1697, or_cse);
  assign nor_802_nl = ~(nor_792_cse | cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6));
  assign mux_1239_nl = MUX_s_1_2_2((mux_1238_nl), (or_2078_nl), nor_802_nl);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl = MUX_v_2_2_2(2'b00, (lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt[7:6]),
      FpNormalize_8U_49U_oelse_not_15);
  assign mux_1240_nl = MUX_s_1_2_2(reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse, IsNaN_8U_23U_4_land_lpi_1_dfm_4,
      reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_8_nl = MUX_v_6_2_2(6'b000000,
      (lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt[5:0]), FpNormalize_8U_49U_oelse_not_15);
  assign FpAdd_8U_23U_o_expo_or_nl = FpAdd_8U_23U_and_57_ssc | (~ mux_1126_cse);
  assign or_1995_nl = (reg_cfg_precision_1_sva_st_13_cse_1[0]) | (~((reg_cfg_precision_1_sva_st_13_cse_1[1])
      & or_tmp_1705));
  assign mux_1242_nl = MUX_s_1_2_2(or_tmp_1707, (~ or_tmp_1705), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_1243_nl = MUX_s_1_2_2((mux_1242_nl), or_tmp_1707, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign mux_1244_nl = MUX_s_1_2_2((mux_1243_nl), (or_1995_nl), lut_lookup_4_if_else_else_acc_itm_10);
  assign and_858_nl = reg_cfg_lut_le_function_1_sva_st_20_cse & IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign mux_198_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, and_858_nl);
  assign and_859_nl = cfg_lut_le_function_1_sva_st_41 & FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign mux_199_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, and_859_nl);
  assign mux_200_nl = MUX_s_1_2_2((mux_199_nl), (mux_198_nl), or_cse);
  assign nor_732_nl = ~(nor_54_cse | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10)
      | reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse | IsNaN_8U_23U_7_land_lpi_1_dfm_6
      | IsNaN_8U_23U_8_land_lpi_1_dfm_4);
  assign nor_733_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_70!=2'b10) |
      IsNaN_8U_23U_7_land_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_lpi_1_dfm_5 | IsNaN_8U_23U_7_land_lpi_1_dfm_st_6
      | FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5);
  assign mux_202_nl = MUX_s_1_2_2((nor_733_nl), (nor_732_nl), or_cse);
  assign nor_729_nl = ~(IsNaN_8U_23U_7_land_lpi_1_dfm_6 | nor_54_cse | reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse
      | IsNaN_8U_23U_8_land_lpi_1_dfm_4 | (~ main_stage_v_2));
  assign mux_203_nl = MUX_s_1_2_2(nor_tmp_55, (nor_729_nl), reg_cfg_precision_1_sva_st_13_cse_1[1]);
  assign mux_204_nl = MUX_s_1_2_2((mux_203_nl), nor_tmp_55, reg_cfg_precision_1_sva_st_13_cse_1[0]);
  assign nor_730_nl = ~(IsNaN_8U_23U_7_land_lpi_1_dfm_7 | IsNaN_8U_23U_8_land_lpi_1_dfm_5
      | IsNaN_8U_23U_7_land_lpi_1_dfm_st_6 | FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5);
  assign mux_205_nl = MUX_s_1_2_2(nor_tmp_57, (nor_730_nl), cfg_precision_1_sva_st_70[1]);
  assign mux_206_nl = MUX_s_1_2_2((mux_205_nl), nor_tmp_57, cfg_precision_1_sva_st_70[0]);
  assign and_59_nl = main_stage_v_3 & (mux_206_nl);
  assign mux_207_nl = MUX_s_1_2_2((and_59_nl), (mux_204_nl), or_cse);
  assign nl_lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl = FpAdd_8U_23U_2_qr_lpi_1_dfm_5
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19)})
      + 8'b1;
  assign lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl = nl_lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_6_nl = MUX_v_8_2_2(8'b00000000,
      (lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl), FpNormalize_8U_49U_2_oelse_not_15);
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_lpi_1_dfm_5
      + 8'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl = nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0];
  assign nand_76_nl = ~(lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp & main_stage_v_2
      & (reg_cfg_precision_1_sva_st_13_cse_1==2'b10));
  assign mux_209_nl = MUX_s_1_2_2(mux_tmp_207, (nand_76_nl), or_cse);
  assign or_306_nl = (~((~(IsNaN_8U_23U_7_land_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_lpi_1_dfm_4))
      | lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp)) | (~ main_stage_v_2) | (reg_cfg_precision_1_sva_st_13_cse_1!=2'b10);
  assign mux_210_nl = MUX_s_1_2_2(mux_tmp_207, (or_306_nl), or_cse);
  assign mux_211_nl = MUX_s_1_2_2((mux_210_nl), (mux_209_nl), nor_54_cse);
  assign mux_213_nl = MUX_s_1_2_2((~ or_1689_cse), main_stage_v_2, IsNaN_8U_23U_7_land_lpi_1_dfm_6);
  assign mux_214_nl = MUX_s_1_2_2((~ or_tmp_63), main_stage_v_3, FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5);
  assign mux_215_nl = MUX_s_1_2_2((mux_214_nl), (mux_213_nl), or_cse);
  assign or_311_nl = (~ lut_lookup_1_if_else_else_else_if_acc_itm_3) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | (~ and_tmp_5);
  assign mux_216_nl = MUX_s_1_2_2((or_311_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign or_315_nl = (~ lut_lookup_else_else_else_asn_mdf_1_sva_st_3) | lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3
      | not_tmp_209;
  assign mux_217_nl = MUX_s_1_2_2((or_315_nl), or_312_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_218_nl = MUX_s_1_2_2((mux_217_nl), (mux_216_nl), or_cse);
  assign nor_726_nl = ~(cfg_lut_le_function_1_sva_st_41 | (~ and_tmp_5));
  assign nor_727_nl = ~(cfg_lut_le_function_1_sva_st_42 | not_tmp_209);
  assign mux_219_nl = MUX_s_1_2_2((nor_727_nl), (nor_726_nl), or_cse);
  assign nor_881_nl = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (~ and_tmp_5));
  assign mux_223_nl = MUX_s_1_2_2((nor_881_nl), and_tmp_5, cfg_lut_le_function_1_sva_st_41);
  assign and_62_nl = IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 & main_stage_v_4 & or_tmp_314;
  assign nor_721_nl = ~(lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 | not_tmp_209);
  assign mux_224_nl = MUX_s_1_2_2((nor_721_nl), (and_62_nl), cfg_lut_le_function_1_sva_st_42);
  assign mux_225_nl = MUX_s_1_2_2((mux_224_nl), (mux_223_nl), or_cse);
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 
      = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp + 8'b10000001;
  assign and_63_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 & main_stage_v_3 & or_1857_cse;
  assign and_64_nl = IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 & main_stage_v_4 & or_tmp_314;
  assign mux_228_nl = MUX_s_1_2_2((and_64_nl), (and_63_nl), or_cse);
  assign or_341_nl = (~ lut_lookup_2_if_else_else_else_if_acc_itm_3_1) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | (~ and_tmp_27);
  assign mux_229_nl = MUX_s_1_2_2((or_341_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign or_346_nl = (~ lut_lookup_else_else_else_asn_mdf_2_sva_st_3) | lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3
      | not_tmp_222;
  assign mux_230_nl = MUX_s_1_2_2((or_346_nl), or_312_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_231_nl = MUX_s_1_2_2((mux_230_nl), (mux_229_nl), or_cse);
  assign nor_719_nl = ~(cfg_lut_le_function_1_sva_st_41 | (~ and_tmp_27));
  assign nor_720_nl = ~(cfg_lut_le_function_1_sva_st_42 | not_tmp_222);
  assign mux_232_nl = MUX_s_1_2_2((nor_720_nl), (nor_719_nl), or_cse);
  assign nor_713_nl = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (~ and_tmp_27));
  assign mux_235_nl = MUX_s_1_2_2((nor_713_nl), and_tmp_27, cfg_lut_le_function_1_sva_st_41);
  assign and_69_nl = IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 & main_stage_v_4 & or_tmp_314;
  assign nor_714_nl = ~(lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3 | not_tmp_222);
  assign mux_236_nl = MUX_s_1_2_2((nor_714_nl), (and_69_nl), cfg_lut_le_function_1_sva_st_42);
  assign mux_237_nl = MUX_s_1_2_2((mux_236_nl), (mux_235_nl), or_cse);
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 
      = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp + 8'b10000001;
  assign and_70_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 & or_1857_cse & main_stage_v_3;
  assign and_71_nl = IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 & main_stage_v_4 & or_tmp_314;
  assign mux_240_nl = MUX_s_1_2_2((and_71_nl), (and_70_nl), or_cse);
  assign or_374_nl = (~ lut_lookup_3_if_else_else_else_if_acc_itm_3_1) | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | (~ and_tmp_14);
  assign mux_241_nl = MUX_s_1_2_2((or_374_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign mux_242_nl = MUX_s_1_2_2(or_tmp_378, or_312_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_243_nl = MUX_s_1_2_2(or_tmp_380, (mux_242_nl), lut_lookup_else_else_else_asn_mdf_3_sva_st_3);
  assign mux_244_nl = MUX_s_1_2_2((mux_243_nl), (mux_241_nl), or_cse);
  assign nor_711_nl = ~(cfg_lut_le_function_1_sva_st_41 | (~ and_tmp_14));
  assign nor_712_nl = ~(cfg_lut_le_function_1_sva_st_42 | not_tmp_235);
  assign mux_245_nl = MUX_s_1_2_2((nor_712_nl), (nor_711_nl), or_cse);
  assign nor_880_nl = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (~ and_tmp_14));
  assign mux_248_nl = MUX_s_1_2_2((nor_880_nl), and_tmp_14, cfg_lut_le_function_1_sva_st_41);
  assign and_74_nl = IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 & main_stage_v_4 & or_tmp_314;
  assign mux_249_nl = MUX_s_1_2_2((~ or_tmp_378), (and_74_nl), cfg_lut_le_function_1_sva_st_42);
  assign mux_250_nl = MUX_s_1_2_2((mux_249_nl), (mux_248_nl), or_cse);
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 
      = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp + 8'b10000001;
  assign and_75_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 & and_tmp_6;
  assign and_76_nl = IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 & main_stage_v_4 & or_tmp_314;
  assign mux_253_nl = MUX_s_1_2_2((and_76_nl), (and_75_nl), or_cse);
  assign or_406_nl = (~ lut_lookup_4_if_else_else_else_if_acc_itm_3_1) | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | (~ and_tmp_19);
  assign mux_254_nl = MUX_s_1_2_2((or_406_nl), or_tmp_63, cfg_lut_le_function_1_sva_st_41);
  assign or_411_nl = (~ lut_lookup_else_else_else_asn_mdf_sva_st_3) | lut_lookup_if_else_else_slc_10_mdf_sva_st_3
      | not_tmp_248;
  assign mux_255_nl = MUX_s_1_2_2((or_411_nl), or_312_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_256_nl = MUX_s_1_2_2((mux_255_nl), (mux_254_nl), or_cse);
  assign nor_705_nl = ~(cfg_lut_le_function_1_sva_st_41 | (~ and_tmp_19));
  assign nor_706_nl = ~(cfg_lut_le_function_1_sva_st_42 | not_tmp_248);
  assign mux_257_nl = MUX_s_1_2_2((nor_706_nl), (nor_705_nl), or_cse);
  assign nor_879_nl = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (~ and_tmp_19));
  assign mux_260_nl = MUX_s_1_2_2((nor_879_nl), and_tmp_19, cfg_lut_le_function_1_sva_st_41);
  assign and_79_nl = IsNaN_8U_23U_6_land_lpi_1_dfm_6 & main_stage_v_4 & or_tmp_314;
  assign nor_700_nl = ~(lut_lookup_if_else_else_slc_10_mdf_sva_st_3 | not_tmp_248);
  assign mux_261_nl = MUX_s_1_2_2((nor_700_nl), (and_79_nl), cfg_lut_le_function_1_sva_st_42);
  assign mux_262_nl = MUX_s_1_2_2((mux_261_nl), (mux_260_nl), or_cse);
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 
      = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp + 8'b10000001;
  assign and_80_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 & and_tmp_6;
  assign and_81_nl = IsNaN_8U_23U_10_land_lpi_1_dfm_5 & main_stage_v_4 & or_tmp_314;
  assign mux_265_nl = MUX_s_1_2_2((and_81_nl), (and_80_nl), or_cse);
  assign lut_lookup_if_else_else_else_else_mux_nl = MUX_v_35_2_2(lut_lookup_1_if_else_else_else_else_else_rshift_itm,
      lut_lookup_1_if_else_else_else_else_if_lshift_itm, IsNaN_8U_23U_6_land_1_lpi_1_dfm_6);
  assign lut_lookup_if_else_else_else_else_mux_1_nl = MUX_v_35_2_2(lut_lookup_2_if_else_else_else_else_else_rshift_itm,
      lut_lookup_2_if_else_else_else_else_if_lshift_itm, IsNaN_8U_23U_6_land_2_lpi_1_dfm_6);
  assign lut_lookup_if_else_else_else_else_mux_2_nl = MUX_v_35_2_2(lut_lookup_3_if_else_else_else_else_else_rshift_itm,
      lut_lookup_3_if_else_else_else_else_if_lshift_itm, IsNaN_8U_23U_6_land_3_lpi_1_dfm_6);
  assign lut_lookup_if_else_else_else_else_mux_3_nl = MUX_v_35_2_2(lut_lookup_4_if_else_else_else_else_else_rshift_itm,
      lut_lookup_4_if_else_else_else_else_if_lshift_itm, IsNaN_8U_23U_6_land_lpi_1_dfm_6);
  assign mux_1138_nl = MUX_s_1_2_2((~ mux_tmp_1136), or_tmp_1513, cfg_lut_uflow_priority_1_sva_9);
  assign and_447_nl = cfg_lut_uflow_priority_1_sva_9 & lut_lookup_lo_uflow_1_lpi_1_dfm_3
      & mux_tmp_1130;
  assign mux_1139_nl = MUX_s_1_2_2((and_447_nl), (mux_1138_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign nor_698_nl = ~((~ (lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9]))
      | lut_lookup_else_if_lor_5_lpi_1_dfm_5 | (~ cfg_lut_le_function_1_sva_st_42)
      | IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 | lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_699_nl = ~(IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 | (~ lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2)
      | lut_lookup_else_if_lor_5_lpi_1_dfm_6 | lut_lookup_else_if_lor_5_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse));
  assign mux_267_nl = MUX_s_1_2_2((nor_699_nl), (nor_698_nl), or_cse);
  assign nor_696_nl = ~(lut_lookup_else_if_lor_5_lpi_1_dfm_5 | (~ cfg_lut_le_function_1_sva_st_42)
      | lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_697_nl = ~(lut_lookup_else_if_lor_5_lpi_1_dfm_6 | lut_lookup_else_if_lor_5_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse));
  assign mux_268_nl = MUX_s_1_2_2((nor_697_nl), (nor_696_nl), or_cse);
  assign or_445_nl = and_854_cse | (~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_269_nl = MUX_s_1_2_2(or_tmp_447, (or_445_nl), or_cse);
  assign nor_694_nl = ~(and_854_cse | (~ cfg_lut_le_function_1_sva_st_42) | IsNaN_8U_23U_6_land_1_lpi_1_dfm_6
      | lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_695_nl = ~(IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 | or_tmp_447);
  assign mux_270_nl = MUX_s_1_2_2((nor_695_nl), (nor_694_nl), or_cse);
  assign mux_272_nl = MUX_s_1_2_2(or_tmp_456, (~ main_stage_v_5), cfg_lut_le_function_1_sva_10);
  assign mux_273_nl = MUX_s_1_2_2((mux_272_nl), or_tmp_456, lut_lookup_unequal_tmp_13);
  assign mux_274_nl = MUX_s_1_2_2((mux_273_nl), mux_tmp_270, or_cse);
  assign mux_276_nl = MUX_s_1_2_2(and_843_cse, and_852_cse, or_cse);
  assign nor_692_nl = ~((~ (lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9]))
      | IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 | lut_lookup_if_1_lor_5_lpi_1_dfm_4 |
      (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_693_nl = ~((~ lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2)
      | lut_lookup_if_1_lor_5_lpi_1_dfm_5 | IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 |
      lut_lookup_if_1_lor_5_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_107!=2'b10)
      | (~ main_stage_v_5));
  assign mux_277_nl = MUX_s_1_2_2((nor_693_nl), (nor_692_nl), or_cse);
  assign nor_691_nl = ~(lut_lookup_if_1_lor_5_lpi_1_dfm_5 | lut_lookup_if_1_lor_5_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5));
  assign mux_278_nl = MUX_s_1_2_2((nor_691_nl), nor_690_cse, or_cse);
  assign nor_689_nl = ~(and_846_cse | lut_lookup_if_1_lor_5_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_107!=2'b10)
      | (~ main_stage_v_5));
  assign mux_279_nl = MUX_s_1_2_2((nor_689_nl), nor_690_cse, or_cse);
  assign or_475_nl = and_846_cse | IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 | lut_lookup_if_1_lor_5_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5);
  assign mux_281_nl = MUX_s_1_2_2((or_475_nl), mux_tmp_279, or_cse);
  assign mux_1151_nl = MUX_s_1_2_2((~ mux_tmp_1149), or_tmp_1523, cfg_lut_uflow_priority_1_sva_9);
  assign and_451_nl = cfg_lut_uflow_priority_1_sva_9 & lut_lookup_lo_uflow_2_lpi_1_dfm_3
      & mux_tmp_1143;
  assign mux_1152_nl = MUX_s_1_2_2((and_451_nl), (mux_1151_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign nor_686_nl = ~((~ (lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9]))
      | (~ cfg_lut_le_function_1_sva_st_42) | IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 |
      lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | lut_lookup_else_if_lor_6_lpi_1_dfm_5 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_687_nl = ~(IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 | (~ lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2)
      | lut_lookup_else_if_lor_6_lpi_1_dfm_6 | lut_lookup_else_if_lor_6_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72[0]) | not_tmp_276);
  assign mux_286_nl = MUX_s_1_2_2((nor_687_nl), (nor_686_nl), or_cse);
  assign nor_684_nl = ~((~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | lut_lookup_else_if_lor_6_lpi_1_dfm_5 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_685_nl = ~(lut_lookup_else_if_lor_6_lpi_1_dfm_6 | lut_lookup_else_if_lor_6_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72[0]) | not_tmp_276);
  assign mux_287_nl = MUX_s_1_2_2((nor_685_nl), (nor_684_nl), or_cse);
  assign nor_681_nl = ~((~ main_stage_v_4) | (~ cfg_lut_le_function_1_sva_st_42)
      | (cfg_precision_1_sva_st_71!=2'b10) | lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | and_82_cse);
  assign nor_682_nl = ~((~ cfg_lut_le_function_1_sva_10) | lut_lookup_else_unequal_tmp_13
      | (~ main_stage_v_5) | (cfg_precision_1_sva_st_72!=2'b10) | lut_lookup_else_if_lor_6_lpi_1_dfm_st_3);
  assign nor_683_nl = ~((~ main_stage_v_5) | (~ cfg_lut_le_function_1_sva_10) | (cfg_precision_1_sva_st_72!=2'b10)
      | lut_lookup_else_if_lor_6_lpi_1_dfm_st_3);
  assign mux_288_nl = MUX_s_1_2_2((nor_683_nl), (nor_682_nl), lut_lookup_else_if_lor_6_lpi_1_dfm_6);
  assign mux_289_nl = MUX_s_1_2_2((mux_288_nl), (nor_681_nl), or_cse);
  assign nor_678_nl = ~((~ main_stage_v_4) | (~ cfg_lut_le_function_1_sva_st_42)
      | (cfg_precision_1_sva_st_71!=2'b10) | lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 | and_82_cse);
  assign nor_679_nl = ~((~ cfg_lut_le_function_1_sva_10) | lut_lookup_else_unequal_tmp_13
      | (~ main_stage_v_5) | (cfg_precision_1_sva_st_72!=2'b10) | lut_lookup_else_if_lor_6_lpi_1_dfm_st_3
      | IsNaN_8U_23U_6_land_2_lpi_1_dfm_7);
  assign nor_680_nl = ~((~ main_stage_v_5) | (~ cfg_lut_le_function_1_sva_10) | (cfg_precision_1_sva_st_72!=2'b10)
      | lut_lookup_else_if_lor_6_lpi_1_dfm_st_3 | IsNaN_8U_23U_6_land_2_lpi_1_dfm_7);
  assign mux_290_nl = MUX_s_1_2_2((nor_680_nl), (nor_679_nl), lut_lookup_else_if_lor_6_lpi_1_dfm_6);
  assign mux_291_nl = MUX_s_1_2_2((mux_290_nl), (nor_678_nl), or_cse);
  assign mux_294_nl = MUX_s_1_2_2(or_tmp_505, (~ main_stage_v_5), cfg_lut_le_function_1_sva_10);
  assign mux_295_nl = MUX_s_1_2_2((mux_294_nl), or_tmp_505, lut_lookup_else_unequal_tmp_13);
  assign mux_296_nl = MUX_s_1_2_2((mux_295_nl), mux_tmp_292, or_cse);
  assign mux_297_nl = MUX_s_1_2_2(or_tmp_505, or_tmp_380, or_cse);
  assign nor_676_nl = ~((~ (lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9]))
      | IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 | lut_lookup_if_1_lor_6_lpi_1_dfm_4 |
      (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_677_nl = ~(IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 | (~ lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2)
      | lut_lookup_if_1_lor_6_lpi_1_dfm_5 | lut_lookup_if_1_lor_6_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5));
  assign mux_299_nl = MUX_s_1_2_2((nor_677_nl), (nor_676_nl), or_cse);
  assign nor_674_nl = ~(lut_lookup_if_1_lor_6_lpi_1_dfm_4 | (~ main_stage_v_4) |
      (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_675_nl = ~(lut_lookup_if_1_lor_6_lpi_1_dfm_5 | lut_lookup_if_1_lor_6_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5));
  assign mux_300_nl = MUX_s_1_2_2((nor_675_nl), (nor_674_nl), or_cse);
  assign mux_301_nl = MUX_s_1_2_2(or_tmp_522, or_365_cse, or_cse);
  assign or_528_nl = IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 | or_tmp_522;
  assign mux_303_nl = MUX_s_1_2_2((or_528_nl), mux_tmp_301, or_cse);
  assign mux_1164_nl = MUX_s_1_2_2((~ mux_tmp_1162), or_tmp_1534, cfg_lut_uflow_priority_1_sva_9);
  assign and_455_nl = cfg_lut_uflow_priority_1_sva_9 & lut_lookup_lo_uflow_3_lpi_1_dfm_3
      & mux_tmp_1156;
  assign mux_1165_nl = MUX_s_1_2_2((and_455_nl), (mux_1164_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign nor_672_nl = ~((~ (lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9]))
      | lut_lookup_else_if_lor_7_lpi_1_dfm_5 | (~ cfg_lut_le_function_1_sva_st_42)
      | IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 | lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_673_nl = ~(IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 | (~ lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2)
      | lut_lookup_else_if_lor_7_lpi_1_dfm_6 | lut_lookup_else_if_lor_7_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse));
  assign mux_308_nl = MUX_s_1_2_2((nor_673_nl), (nor_672_nl), or_cse);
  assign nor_670_nl = ~(lut_lookup_else_if_lor_7_lpi_1_dfm_5 | (~ cfg_lut_le_function_1_sva_st_42)
      | lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_671_nl = ~(lut_lookup_else_if_lor_7_lpi_1_dfm_6 | lut_lookup_else_if_lor_7_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse));
  assign mux_309_nl = MUX_s_1_2_2((nor_671_nl), (nor_670_nl), or_cse);
  assign or_545_nl = and_839_cse | (~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_310_nl = MUX_s_1_2_2(or_tmp_547, (or_545_nl), or_cse);
  assign nor_668_nl = ~(and_839_cse | (~ cfg_lut_le_function_1_sva_st_42) | IsNaN_8U_23U_6_land_3_lpi_1_dfm_6
      | lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_669_nl = ~(IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 | or_tmp_547);
  assign mux_311_nl = MUX_s_1_2_2((nor_669_nl), (nor_668_nl), or_cse);
  assign nor_666_nl = ~((~ (lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9]))
      | IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 | lut_lookup_if_1_lor_7_lpi_1_dfm_4 |
      (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_667_nl = ~((~ lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2)
      | lut_lookup_if_1_lor_7_lpi_1_dfm_5 | IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 |
      lut_lookup_if_1_lor_7_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_107!=2'b10)
      | (~ main_stage_v_5));
  assign mux_319_nl = MUX_s_1_2_2((nor_667_nl), (nor_666_nl), or_cse);
  assign or_566_nl = lut_lookup_if_1_lor_7_lpi_1_dfm_5 | lut_lookup_if_1_lor_7_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5);
  assign mux_320_nl = MUX_s_1_2_2((or_566_nl), or_tmp_397, or_cse);
  assign or_569_nl = and_850_cse | lut_lookup_if_1_lor_7_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_107!=2'b10)
      | (~ main_stage_v_5);
  assign mux_322_nl = MUX_s_1_2_2((or_569_nl), or_tmp_397, or_cse);
  assign or_575_nl = and_850_cse | IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 | lut_lookup_if_1_lor_7_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5);
  assign mux_325_nl = MUX_s_1_2_2((or_575_nl), or_tmp_573, or_cse);
  assign mux_1177_nl = MUX_s_1_2_2((~ mux_tmp_1175), or_tmp_1545, cfg_lut_uflow_priority_1_sva_9);
  assign and_459_nl = cfg_lut_uflow_priority_1_sva_9 & lut_lookup_lo_uflow_lpi_1_dfm_3
      & mux_tmp_1169;
  assign mux_1178_nl = MUX_s_1_2_2((and_459_nl), (mux_1177_nl), cfg_lut_hybrid_priority_1_sva_9);
  assign nor_664_nl = ~((~ (lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9]))
      | lut_lookup_else_if_lor_1_lpi_1_dfm_5 | (~ cfg_lut_le_function_1_sva_st_42)
      | IsNaN_8U_23U_6_land_lpi_1_dfm_6 | lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_665_nl = ~(IsNaN_8U_23U_6_land_lpi_1_dfm_7 | (~ lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2)
      | lut_lookup_else_if_lor_1_lpi_1_dfm_6 | lut_lookup_else_if_lor_1_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse));
  assign mux_332_nl = MUX_s_1_2_2((nor_665_nl), (nor_664_nl), or_cse);
  assign nor_662_nl = ~(lut_lookup_else_if_lor_1_lpi_1_dfm_5 | (~ cfg_lut_le_function_1_sva_st_42)
      | lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_663_nl = ~(lut_lookup_else_if_lor_1_lpi_1_dfm_6 | lut_lookup_else_if_lor_1_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_72!=2'b10) | (~ and_843_cse));
  assign mux_333_nl = MUX_s_1_2_2((nor_663_nl), (nor_662_nl), or_cse);
  assign or_596_nl = and_835_cse | (~ cfg_lut_le_function_1_sva_st_42) | lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_334_nl = MUX_s_1_2_2(or_tmp_598, (or_596_nl), or_cse);
  assign nor_660_nl = ~(and_835_cse | (~ cfg_lut_le_function_1_sva_st_42) | IsNaN_8U_23U_6_land_lpi_1_dfm_6
      | lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_661_nl = ~(IsNaN_8U_23U_6_land_lpi_1_dfm_7 | or_tmp_598);
  assign mux_335_nl = MUX_s_1_2_2((nor_661_nl), (nor_660_nl), or_cse);
  assign nor_658_nl = ~((~ (lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9]))
      | IsNaN_8U_23U_10_land_lpi_1_dfm_5 | lut_lookup_if_1_lor_1_lpi_1_dfm_4 | (~
      main_stage_v_4) | (cfg_precision_1_sva_st_71!=2'b10));
  assign nor_659_nl = ~((~ lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2)
      | lut_lookup_if_1_lor_1_lpi_1_dfm_5 | IsNaN_8U_23U_10_land_lpi_1_dfm_6 | lut_lookup_if_1_lor_1_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5));
  assign mux_343_nl = MUX_s_1_2_2((nor_659_nl), (nor_658_nl), or_cse);
  assign or_617_nl = lut_lookup_if_1_lor_1_lpi_1_dfm_5 | lut_lookup_if_1_lor_1_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5);
  assign mux_344_nl = MUX_s_1_2_2((or_617_nl), or_tmp_428, or_cse);
  assign or_620_nl = and_848_cse | lut_lookup_if_1_lor_1_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_107!=2'b10)
      | (~ main_stage_v_5);
  assign mux_346_nl = MUX_s_1_2_2((or_620_nl), or_tmp_428, or_cse);
  assign or_625_nl = and_848_cse | IsNaN_8U_23U_10_land_lpi_1_dfm_6 | lut_lookup_if_1_lor_1_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_107!=2'b10) | (~ main_stage_v_5);
  assign mux_349_nl = MUX_s_1_2_2((or_625_nl), or_tmp_623, or_cse);
  assign lut_lookup_else_else_lut_lookup_else_else_and_10_nl = (~ lut_lookup_else_else_else_asn_mdf_sva_4)
      & lut_lookup_else_else_slc_32_mdf_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_11_nl = (~(lut_lookup_if_else_else_else_asn_mdf_sva_2
      | lut_lookup_if_else_else_slc_10_mdf_sva_4)) & lut_lookup_4_if_else_slc_32_svs_8;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_4_nl = ~(lut_lookup_4_if_if_else_else_if_acc_itm_3
      | lut_lookup_4_if_if_else_acc_itm_9_1 | lut_lookup_if_if_lor_1_lpi_1_dfm_4);
  assign lut_lookup_else_else_lut_lookup_else_else_and_7_nl = (~ lut_lookup_else_else_else_asn_mdf_3_sva_4)
      & lut_lookup_else_else_slc_32_mdf_3_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_12_nl = (~(lut_lookup_if_else_else_else_asn_mdf_2_sva_2
      | lut_lookup_if_else_else_slc_10_mdf_2_sva_4)) & lut_lookup_2_if_else_slc_32_svs_8;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_5_nl = ~(lut_lookup_2_if_if_else_else_if_acc_itm_3
      | lut_lookup_2_if_if_else_acc_itm_9_1 | lut_lookup_if_if_lor_6_lpi_1_dfm_4);
  assign lut_lookup_else_else_lut_lookup_else_else_and_4_nl = (~ lut_lookup_else_else_else_asn_mdf_2_sva_4)
      & lut_lookup_else_else_slc_32_mdf_2_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_13_nl = (~(lut_lookup_if_else_else_else_asn_mdf_1_sva_2
      | lut_lookup_if_else_else_slc_10_mdf_1_sva_4)) & lut_lookup_1_if_else_slc_32_svs_8;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_6_nl = ~(lut_lookup_1_if_if_else_else_if_acc_itm_3
      | lut_lookup_1_if_if_else_acc_itm_9_1 | lut_lookup_if_if_lor_5_lpi_1_dfm_4);
  assign lut_lookup_else_else_lut_lookup_else_else_and_1_nl = (~ lut_lookup_else_else_else_asn_mdf_1_sva_4)
      & lut_lookup_else_else_slc_32_mdf_1_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_14_nl = (~(lut_lookup_if_else_else_else_asn_mdf_3_sva_2
      | lut_lookup_if_else_else_slc_10_mdf_3_sva_4)) & lut_lookup_3_if_else_slc_32_svs_8;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_7_nl = ~(lut_lookup_3_if_if_else_else_if_acc_itm_3
      | lut_lookup_3_if_if_else_acc_itm_9_1 | lut_lookup_if_if_lor_7_lpi_1_dfm_4);
  assign and_830_nl = or_1853_cse & main_stage_v_4;
  assign mux_371_nl = MUX_s_1_2_2(not_tmp_334, main_stage_v_5, lut_lookup_unequal_tmp_13);
  assign mux_372_nl = MUX_s_1_2_2((mux_371_nl), (and_830_nl), or_cse);
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_8_nl = MUX_v_8_2_2((cfg_lut_le_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[30:23]), FpAdd_8U_23U_b_right_shift_qif_and_tmp);
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_9_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[30:23])),
      (~ (cfg_lut_le_start_rsci_d[30:23])), FpAdd_8U_23U_b_right_shift_qif_and_tmp);
  assign nl_acc_4_nl = ({(FpAdd_8U_23U_a_right_shift_qelse_mux_8_nl) , 1'b1}) + ({(FpAdd_8U_23U_a_right_shift_qelse_mux_9_nl)
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[8:0];
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_14_nl = MUX_v_8_2_2((cfg_lut_lo_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[62:55]), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3);
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_15_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[62:55])),
      (~ (cfg_lut_lo_start_rsci_d[30:23])), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3);
  assign nl_acc_10_nl = ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_14_nl) , 1'b1})
      + ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_15_nl) , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[8:0];
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_12_nl = MUX_v_8_2_2((cfg_lut_lo_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[94:87]), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2);
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_13_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[94:87])),
      (~ (cfg_lut_lo_start_rsci_d[30:23])), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2);
  assign nl_acc_9_nl = ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_12_nl) , 1'b1})
      + ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_13_nl) , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[8:0];
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_8_nl = MUX_v_8_2_2((cfg_lut_lo_start_rsci_d[30:23]),
      (chn_lut_in_rsci_d_mxwt[126:119]), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp);
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_9_nl = MUX_v_8_2_2((~ (chn_lut_in_rsci_d_mxwt[126:119])),
      (~ (cfg_lut_lo_start_rsci_d[30:23])), FpAdd_8U_23U_2_b_right_shift_qif_and_tmp);
  assign nl_acc_5_nl = ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_8_nl) , 1'b1}) +
      ({(FpAdd_8U_23U_2_a_right_shift_qelse_mux_9_nl) , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[8:0];
  assign or_827_nl = main_stage_v_1 | (~ mux_tmp_595);
  assign mux_598_nl = MUX_s_1_2_2((or_827_nl), main_stage_v_1, nor_648_cse);
  assign mux_599_nl = MUX_s_1_2_2(mux_tmp_596, (~ (mux_598_nl)), reg_cfg_precision_1_sva_st_12_cse_1[1]);
  assign mux_600_nl = MUX_s_1_2_2((mux_599_nl), mux_tmp_596, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign or_829_nl = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign mux_601_nl = MUX_s_1_2_2((~ main_stage_v_2), or_1689_cse, or_829_nl);
  assign mux_602_nl = MUX_s_1_2_2(or_1689_cse, (mux_601_nl), main_stage_v_1);
  assign mux_605_nl = MUX_s_1_2_2(or_1689_cse, (mux_602_nl), nor_190_cse);
  assign mux_606_nl = MUX_s_1_2_2((mux_605_nl), (mux_600_nl), or_cse);
  assign or_839_nl = nor_193_cse | (~(IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_8_land_1_lpi_1_dfm_6))
      | (~ reg_chn_lut_out_rsci_ld_core_psct_cse) | chn_lut_out_rsci_bawt;
  assign mux_611_nl = MUX_s_1_2_2(or_cse, (or_839_nl), main_stage_v_2);
  assign mux_620_nl = MUX_s_1_2_2(mux_tmp_618, (~ (mux_611_nl)), reg_cfg_precision_1_sva_st_12_cse_1[1]);
  assign mux_621_nl = MUX_s_1_2_2((mux_620_nl), mux_tmp_618, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign mux_622_nl = MUX_s_1_2_2(mux_tmp_617, (mux_621_nl), main_stage_v_1);
  assign mux_477_nl = MUX_s_1_2_2(not_tmp_394, mux_tmp_475, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign nand_15_nl = ~(main_stage_v_1 & (~ (mux_477_nl)));
  assign mux_624_nl = MUX_s_1_2_2((nand_15_nl), or_1688_cse, IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4);
  assign mux_625_nl = MUX_s_1_2_2(not_tmp_394, mux_tmp_475, or_849_cse);
  assign mux_627_nl = MUX_s_1_2_2((mux_625_nl), (mux_624_nl), nor_648_cse);
  assign or_850_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 | IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  assign mux_628_nl = MUX_s_1_2_2((~ main_stage_v_2), or_1689_cse, or_850_nl);
  assign mux_631_nl = MUX_s_1_2_2(or_1689_cse, (mux_628_nl), nor_196_cse);
  assign mux_634_nl = MUX_s_1_2_2((mux_631_nl), (mux_627_nl), or_cse);
  assign mux_518_nl = MUX_s_1_2_2((~ not_tmp_412), or_1689_cse, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign nand_16_nl = ~(main_stage_v_1 & (mux_518_nl));
  assign mux_635_nl = MUX_s_1_2_2((nand_16_nl), or_1688_cse, reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse);
  assign mux_636_nl = MUX_s_1_2_2(not_tmp_412, (~ or_1689_cse), or_849_cse);
  assign mux_638_nl = MUX_s_1_2_2((mux_636_nl), (mux_635_nl), nor_648_cse);
  assign mux_645_nl = MUX_s_1_2_2(mux_tmp_643, (mux_638_nl), or_cse);
  assign mux_534_nl = MUX_s_1_2_2(not_tmp_418, or_1689_cse, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign nand_17_nl = ~(main_stage_v_1 & (~ (mux_534_nl)));
  assign mux_646_nl = MUX_s_1_2_2((nand_17_nl), or_1688_cse, reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse);
  assign mux_647_nl = MUX_s_1_2_2(not_tmp_418, or_1689_cse, or_849_cse);
  assign mux_649_nl = MUX_s_1_2_2((mux_647_nl), (mux_646_nl), nor_648_cse);
  assign mux_650_nl = MUX_s_1_2_2(mux_tmp_643, (mux_649_nl), or_cse);
  assign mux_651_nl = MUX_s_1_2_2((mux_650_nl), (mux_645_nl), nor_54_cse);
  assign mux_652_nl = MUX_s_1_2_2(and_tmp_59, main_stage_v_1, or_cse);
  assign nor_642_nl = ~((~ reg_chn_lut_out_rsci_ld_core_psct_cse) | chn_lut_out_rsci_bawt
      | (~ and_tmp_59));
  assign and_827_nl = or_26_cse & reg_cfg_lut_le_function_1_sva_st_19_cse & FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  assign mux_653_nl = MUX_s_1_2_2((nor_642_nl), (mux_652_nl), and_827_nl);
  assign nl_lut_lookup_else_1_lo_index_u_1_sva_3  = (lut_in_data_sva_154[31:0]) -
      cfg_lut_lo_start_1_sva_41;
  assign mux_548_nl = MUX_s_1_2_2(not_tmp_422, main_stage_v_1, reg_cfg_precision_1_sva_st_12_cse_1[0]);
  assign and_98_nl = FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 & (mux_548_nl);
  assign mux_654_nl = MUX_s_1_2_2(and_tmp_61, (and_98_nl), or_cse);
  assign and_100_nl = reg_cfg_lut_le_function_1_sva_st_19_cse & FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5
      & or_26_cse & main_stage_v_1;
  assign and_101_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & reg_cfg_lut_le_function_1_sva_st_20_cse
      & main_stage_v_2 & or_66_cse;
  assign mux_655_nl = MUX_s_1_2_2((and_101_nl), (and_100_nl), or_cse);
  assign nl_lut_lookup_else_1_lo_index_u_2_sva_3  = (lut_in_data_sva_154[63:32])
      - cfg_lut_lo_start_1_sva_41;
  assign and_102_nl = FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 & main_stage_v_1
      & or_26_cse;
  assign and_103_nl = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 & mux_tmp_655;
  assign mux_657_nl = MUX_s_1_2_2((and_103_nl), (and_102_nl), or_cse);
  assign and_104_nl = main_stage_v_1 & FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5
      & reg_cfg_lut_le_function_1_sva_st_19_cse & or_26_cse;
  assign and_105_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & reg_cfg_lut_le_function_1_sva_st_20_cse
      & main_stage_v_2 & or_66_cse;
  assign mux_658_nl = MUX_s_1_2_2((and_105_nl), (and_104_nl), or_cse);
  assign nl_lut_lookup_else_1_lo_index_u_3_sva_3  = (lut_in_data_sva_154[95:64])
      - cfg_lut_lo_start_1_sva_41;
  assign and_106_nl = FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 & main_stage_v_1
      & or_26_cse;
  assign mux_659_nl = MUX_s_1_2_2(and_tmp_69, (and_106_nl), or_cse);
  assign and_108_nl = main_stage_v_1 & FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5
      & reg_cfg_lut_le_function_1_sva_st_19_cse & or_26_cse;
  assign and_109_nl = reg_cfg_lut_le_function_1_sva_st_20_cse & IsNaN_8U_23U_1_land_lpi_1_dfm_7
      & main_stage_v_2 & or_66_cse;
  assign mux_660_nl = MUX_s_1_2_2((and_109_nl), (and_108_nl), or_cse);
  assign nl_lut_lookup_else_1_lo_index_u_sva_3  = (lut_in_data_sva_154[127:96]) -
      cfg_lut_lo_start_1_sva_41;
  assign and_110_nl = FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 & main_stage_v_1
      & or_26_cse;
  assign and_111_nl = IsNaN_8U_23U_7_land_lpi_1_dfm_6 & main_stage_v_2 & or_66_cse;
  assign mux_661_nl = MUX_s_1_2_2((and_111_nl), (and_110_nl), or_cse);
  assign or_879_nl = (~(IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp | FpAdd_8U_23U_1_mux_61_itm_4
      | IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp)) | (cfg_precision_1_sva_st_70!=2'b10);
  assign nor_638_nl = ~(lut_lookup_4_if_else_slc_32_svs_7 | (~ or_1857_cse));
  assign or_880_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (~ lut_lookup_4_if_else_else_else_if_acc_itm_3_1)
      | (~ FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6) | lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign mux_662_nl = MUX_s_1_2_2((nor_638_nl), or_1857_cse, or_880_nl);
  assign mux_663_nl = MUX_s_1_2_2((~ (mux_662_nl)), (or_879_nl), cfg_lut_le_function_1_sva_st_41);
  assign and_112_nl = main_stage_v_3 & (mux_663_nl);
  assign or_885_nl = (~(lut_lookup_else_unequal_tmp_12 | lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2))
      | (cfg_precision_1_sva_st_71!=2'b10);
  assign or_887_nl = (~ lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2)
      | (cfg_precision_1_sva_st_71!=2'b10);
  assign mux_664_nl = MUX_s_1_2_2((or_887_nl), (or_885_nl), lut_lookup_else_if_lor_1_lpi_1_dfm_5);
  assign nor_640_nl = ~(lut_lookup_4_if_else_slc_32_svs_8 | (~ or_tmp_314));
  assign or_888_nl = (~ lut_lookup_4_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_sva_st_3
      | (~ lut_lookup_if_else_else_else_asn_mdf_sva_2) | lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign mux_665_nl = MUX_s_1_2_2((nor_640_nl), or_tmp_314, or_888_nl);
  assign mux_666_nl = MUX_s_1_2_2((~ (mux_665_nl)), (mux_664_nl), cfg_lut_le_function_1_sva_st_42);
  assign and_113_nl = main_stage_v_4 & (mux_666_nl);
  assign mux_667_nl = MUX_s_1_2_2((and_113_nl), (and_112_nl), or_cse);
  assign mux_672_nl = MUX_s_1_2_2(main_stage_v_4, and_826_cse, or_cse);
  assign or_899_nl = (~(IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp | FpAdd_8U_23U_1_mux_45_itm_4
      | IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp)) | (cfg_precision_1_sva_st_70!=2'b10);
  assign nor_633_nl = ~(lut_lookup_3_if_else_slc_32_svs_7 | (~ or_1857_cse));
  assign or_900_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (~ lut_lookup_3_if_else_else_else_if_acc_itm_3_1)
      | (~ FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6) | lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign mux_673_nl = MUX_s_1_2_2((nor_633_nl), or_1857_cse, or_900_nl);
  assign mux_674_nl = MUX_s_1_2_2((~ (mux_673_nl)), (or_899_nl), cfg_lut_le_function_1_sva_st_41);
  assign and_114_nl = main_stage_v_3 & (mux_674_nl);
  assign nand_18_nl = ~(lut_lookup_else_if_lor_7_lpi_1_dfm_5 & nor_634_cse);
  assign mux_675_nl = MUX_s_1_2_2((nand_18_nl), or_tmp_314, lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2);
  assign nor_636_nl = ~(lut_lookup_3_if_else_slc_32_svs_8 | (~ or_tmp_314));
  assign or_907_nl = (~ lut_lookup_3_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3
      | (~ lut_lookup_if_else_else_else_asn_mdf_3_sva_2) | lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign mux_676_nl = MUX_s_1_2_2((nor_636_nl), or_tmp_314, or_907_nl);
  assign mux_677_nl = MUX_s_1_2_2((~ (mux_676_nl)), (mux_675_nl), cfg_lut_le_function_1_sva_st_42);
  assign and_115_nl = main_stage_v_4 & (mux_677_nl);
  assign mux_678_nl = MUX_s_1_2_2((and_115_nl), (and_114_nl), or_cse);
  assign or_915_nl = (~(IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp | FpAdd_8U_23U_1_mux_29_itm_4
      | IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp)) | (cfg_precision_1_sva_st_70!=2'b10);
  assign nor_628_nl = ~(lut_lookup_2_if_else_slc_32_svs_7 | (~ or_1857_cse));
  assign or_916_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (~ lut_lookup_2_if_else_else_else_if_acc_itm_3_1)
      | (~ FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6) | lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign mux_684_nl = MUX_s_1_2_2((nor_628_nl), or_1857_cse, or_916_nl);
  assign mux_685_nl = MUX_s_1_2_2((~ (mux_684_nl)), (or_915_nl), cfg_lut_le_function_1_sva_st_41);
  assign and_116_nl = main_stage_v_3 & (mux_685_nl);
  assign nand_19_nl = ~(lut_lookup_else_if_lor_6_lpi_1_dfm_5 & nor_634_cse);
  assign mux_686_nl = MUX_s_1_2_2((nand_19_nl), or_tmp_314, lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2);
  assign nor_631_nl = ~(lut_lookup_2_if_else_slc_32_svs_8 | (~ or_tmp_314));
  assign or_923_nl = (~ lut_lookup_2_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3
      | (~ lut_lookup_if_else_else_else_asn_mdf_2_sva_2) | lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign mux_687_nl = MUX_s_1_2_2((nor_631_nl), or_tmp_314, or_923_nl);
  assign mux_688_nl = MUX_s_1_2_2((~ (mux_687_nl)), (mux_686_nl), cfg_lut_le_function_1_sva_st_42);
  assign and_117_nl = main_stage_v_4 & (mux_688_nl);
  assign mux_689_nl = MUX_s_1_2_2((and_117_nl), (and_116_nl), or_cse);
  assign or_931_nl = (~ lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1) | (cfg_precision_1_sva_st_70!=2'b10);
  assign nor_623_nl = ~(lut_lookup_1_if_else_slc_32_svs_7 | (~ or_1857_cse));
  assign or_932_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (~ lut_lookup_1_if_else_else_else_if_acc_itm_3)
      | (~ FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6) | lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign mux_695_nl = MUX_s_1_2_2((nor_623_nl), or_1857_cse, or_932_nl);
  assign mux_696_nl = MUX_s_1_2_2((~ (mux_695_nl)), (or_931_nl), cfg_lut_le_function_1_sva_st_41);
  assign and_118_nl = main_stage_v_3 & (mux_696_nl);
  assign nand_20_nl = ~(lut_lookup_else_if_lor_5_lpi_1_dfm_5 & (~((~ lut_lookup_else_unequal_tmp_18)
      | (cfg_precision_1_sva_st_71!=2'b10))));
  assign mux_697_nl = MUX_s_1_2_2((nand_20_nl), or_tmp_314, lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2);
  assign nor_626_nl = ~(lut_lookup_1_if_else_slc_32_svs_8 | (~ or_tmp_314));
  assign or_939_nl = (~ lut_lookup_1_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3
      | (~ lut_lookup_if_else_else_else_asn_mdf_1_sva_2) | lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign mux_698_nl = MUX_s_1_2_2((nor_626_nl), or_tmp_314, or_939_nl);
  assign mux_699_nl = MUX_s_1_2_2((~ (mux_698_nl)), (mux_697_nl), cfg_lut_le_function_1_sva_st_42);
  assign and_119_nl = main_stage_v_4 & (mux_699_nl);
  assign mux_700_nl = MUX_s_1_2_2((and_119_nl), (and_118_nl), or_cse);
  assign mux_704_nl = MUX_s_1_2_2(mux_tmp_270, mux_670_cse, or_cse);
  assign and_823_nl = ((~(FpAdd_8U_23U_2_mux_61_itm_3 | and_1138_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp))
      | (cfg_precision_1_sva_st_70!=2'b10)) & main_stage_v_3;
  assign mux_710_nl = MUX_s_1_2_2(main_stage_v_4, and_tmp_83, lut_lookup_if_1_lor_1_lpi_1_dfm_4);
  assign mux_711_nl = MUX_s_1_2_2((mux_710_nl), (and_823_nl), or_cse);
  assign and_822_nl = ((~(FpAdd_8U_23U_2_mux_45_itm_3 | and_1139_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp))
      | (cfg_precision_1_sva_st_70!=2'b10)) & main_stage_v_3;
  assign mux_721_nl = MUX_s_1_2_2(main_stage_v_4, and_tmp_83, lut_lookup_if_1_lor_7_lpi_1_dfm_4);
  assign mux_722_nl = MUX_s_1_2_2((mux_721_nl), (and_822_nl), or_cse);
  assign nor_619_nl = ~(and_1140_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp
      | FpAdd_8U_23U_2_mux_29_itm_3 | (~ main_stage_v_3));
  assign mux_730_nl = MUX_s_1_2_2((nor_619_nl), main_stage_v_3, or_1857_cse);
  assign mux_731_nl = MUX_s_1_2_2(main_stage_v_4, and_tmp_83, lut_lookup_if_1_lor_6_lpi_1_dfm_4);
  assign mux_732_nl = MUX_s_1_2_2((mux_731_nl), (mux_730_nl), or_cse);
  assign mux_737_nl = MUX_s_1_2_2(main_stage_v_3, and_tmp_6, or_969_cse);
  assign mux_738_nl = MUX_s_1_2_2(main_stage_v_4, and_tmp_83, lut_lookup_if_1_lor_5_lpi_1_dfm_4);
  assign mux_739_nl = MUX_s_1_2_2((mux_738_nl), (mux_737_nl), or_cse);
  assign nor_616_nl = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (~ FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6)
      | lut_lookup_if_else_else_slc_10_mdf_1_sva_3 | (~(lut_lookup_1_if_else_slc_32_svs_7
      & mux_tmp_704)));
  assign mux_751_nl = MUX_s_1_2_2((nor_616_nl), main_stage_v_3, or_1857_cse);
  assign and_1166_nl = (mux_751_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign mux_756_nl = MUX_s_1_2_2(or_tmp_993, (~ mux_755_cse), lut_lookup_1_if_else_slc_32_svs_8);
  assign or_990_nl = (~ lut_lookup_1_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3
      | lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign mux_757_nl = MUX_s_1_2_2((mux_756_nl), or_tmp_993, or_990_nl);
  assign mux_758_nl = MUX_s_1_2_2((mux_757_nl), or_978_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_759_nl = MUX_s_1_2_2((~ (mux_758_nl)), (and_1166_nl), or_cse);
  assign and_127_nl = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & lut_lookup_1_if_else_slc_32_svs_7
      & mux_tmp_704;
  assign mux_761_nl = MUX_s_1_2_2((and_127_nl), main_stage_v_3, or_1857_cse);
  assign and_1164_nl = (mux_761_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign and_819_nl = lut_lookup_1_if_else_slc_32_svs_st_5 & lut_lookup_1_if_else_slc_32_svs_8;
  assign mux_766_nl = MUX_s_1_2_2((~ or_tmp_993), mux_755_cse, and_819_nl);
  assign mux_767_nl = MUX_s_1_2_2((mux_766_nl), nor_612_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_768_nl = MUX_s_1_2_2((mux_767_nl), (and_1164_nl), or_cse);
  assign mux_1245_nl = MUX_s_1_2_2(nor_832_cse, and_1142_cse, cfg_lut_le_function_1_sva_st_41);
  assign nor_831_nl = ~(IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp | FpAdd_8U_23U_1_mux_13_itm_4
      | (mux_1245_nl));
  assign nor_833_nl = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (~ lut_lookup_1_if_else_else_else_if_acc_itm_3)
      | (~ FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6) | lut_lookup_if_else_else_slc_10_mdf_1_sva_3
      | (~ lut_lookup_1_if_else_slc_32_svs_7) | cfg_lut_le_function_1_sva_st_41);
  assign mux_1246_nl = MUX_s_1_2_2((nor_833_nl), (nor_831_nl), nor_792_cse);
  assign nor_597_nl = ~((~ lut_lookup_1_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | (~ lut_lookup_1_if_else_else_else_if_acc_itm_3) | (~ lut_lookup_1_if_else_slc_32_svs_7)
      | lut_lookup_if_else_else_slc_10_mdf_1_sva_3 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | (~ and_tmp_5));
  assign nor_598_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~ IsNaN_8U_23U_6_land_1_lpi_1_dfm_6)
      | (~ lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2)
      | (~ lut_lookup_else_else_else_asn_mdf_1_sva_st_3) | (~ lut_lookup_if_else_else_else_asn_mdf_1_sva_2)
      | lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 | lut_lookup_if_else_else_slc_10_mdf_1_sva_4
      | (~(lut_lookup_1_if_else_slc_32_svs_8 & lut_lookup_1_if_else_slc_32_svs_st_5
      & main_stage_v_4 & or_tmp_314)));
  assign mux_783_nl = MUX_s_1_2_2((nor_598_nl), (nor_597_nl), or_cse);
  assign and_815_nl = (~ cfg_lut_le_function_1_sva_st_41) & main_stage_v_3;
  assign and_816_nl = (~ cfg_lut_le_function_1_sva_st_42) & main_stage_v_4;
  assign mux_784_nl = MUX_s_1_2_2((and_816_nl), (and_815_nl), or_cse);
  assign and_131_nl = lut_lookup_else_else_else_asn_mdf_1_sva_4 & lut_lookup_else_else_slc_32_mdf_1_sva_8
      & cfg_lut_le_function_1_sva_st_42 & IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 & lut_lookup_else_else_else_asn_mdf_1_sva_st_3
      & main_stage_v_4 & or_tmp_314;
  assign mux_785_nl = MUX_s_1_2_2((and_131_nl), and_tmp_92, or_cse);
  assign nor_595_nl = ~((cfg_precision_1_sva_st_71[1]) | (~ nor_tmp_238));
  assign mux_790_nl = MUX_s_1_2_2((nor_595_nl), nor_tmp_238, cfg_precision_1_sva_st_71[0]);
  assign mux_791_nl = MUX_s_1_2_2((mux_790_nl), main_stage_v_4, and_814_cse);
  assign mux_792_nl = MUX_s_1_2_2((mux_791_nl), mux_789_cse, or_cse);
  assign mux_796_nl = MUX_s_1_2_2(and_134_cse, main_stage_v_4, and_814_cse);
  assign mux_797_nl = MUX_s_1_2_2((mux_796_nl), mux_851_cse, or_cse);
  assign mux_798_nl = MUX_s_1_2_2(mux_tmp_279, or_tmp_331, or_cse);
  assign or_1045_nl = lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
      | lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
      | (~ and_tmp_98);
  assign mux_799_nl = MUX_s_1_2_2((or_1045_nl), or_tmp_1043, or_cse);
  assign or_2009_nl = nor_792_cse | (~ FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_1_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_1_sva_7);
  assign nor_830_nl = ~((cfg_precision_1_sva_st_70[1]) | (~ or_tmp_1716));
  assign mux_1247_nl = MUX_s_1_2_2((nor_830_nl), or_tmp_1716, cfg_precision_1_sva_st_70[0]);
  assign or_2007_nl = and_1141_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp;
  assign mux_1248_nl = MUX_s_1_2_2((mux_1247_nl), (or_2009_nl), or_2007_nl);
  assign mux_803_nl = MUX_s_1_2_2(and_tmp_98, and_tmp_97, or_cse);
  assign mux_806_nl = MUX_s_1_2_2(mux_805_cse, mux_793_cse, or_cse);
  assign mux_815_nl = MUX_s_1_2_2(nor_588_cse, main_stage_v_3, or_1857_cse);
  assign and_1162_nl = (mux_815_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign mux_820_nl = MUX_s_1_2_2(or_tmp_993, (~ mux_755_cse), lut_lookup_2_if_else_slc_32_svs_8);
  assign or_1072_nl = (~ lut_lookup_2_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3
      | lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign mux_821_nl = MUX_s_1_2_2((mux_820_nl), or_tmp_993, or_1072_nl);
  assign mux_822_nl = MUX_s_1_2_2((mux_821_nl), or_978_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_823_nl = MUX_s_1_2_2((~ (mux_822_nl)), (and_1162_nl), or_cse);
  assign and_138_nl = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & lut_lookup_2_if_else_slc_32_svs_7
      & mux_tmp_704;
  assign mux_825_nl = MUX_s_1_2_2((and_138_nl), main_stage_v_3, or_1857_cse);
  assign and_1160_nl = (mux_825_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign and_812_nl = lut_lookup_2_if_else_slc_32_svs_st_5 & lut_lookup_2_if_else_slc_32_svs_8;
  assign mux_830_nl = MUX_s_1_2_2((~ or_tmp_993), mux_755_cse, and_812_nl);
  assign mux_831_nl = MUX_s_1_2_2((mux_830_nl), nor_612_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_832_nl = MUX_s_1_2_2((mux_831_nl), (and_1160_nl), or_cse);
  assign nor_575_nl = ~((~ lut_lookup_2_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | (~ lut_lookup_2_if_else_else_else_if_acc_itm_3_1) | lut_lookup_if_else_else_slc_10_mdf_2_sva_3
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (~(lut_lookup_2_if_else_slc_32_svs_7
      & FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & main_stage_v_3 & or_1857_cse)));
  assign nor_576_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~ lut_lookup_if_else_else_else_asn_mdf_2_sva_2)
      | (~ lut_lookup_else_else_else_asn_mdf_2_sva_st_3) | lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3
      | lut_lookup_if_else_else_slc_10_mdf_2_sva_4 | (~(lut_lookup_2_if_else_slc_32_svs_8
      & IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 & lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      & lut_lookup_2_if_else_slc_32_svs_st_5 & main_stage_v_4 & or_tmp_314)));
  assign mux_840_nl = MUX_s_1_2_2((nor_576_nl), (nor_575_nl), or_cse);
  assign and_142_nl = lut_lookup_else_else_else_asn_mdf_2_sva_4 & cfg_lut_le_function_1_sva_st_42
      & lut_lookup_else_else_else_asn_mdf_2_sva_st_3 & lut_lookup_else_else_slc_32_mdf_2_sva_8
      & IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 & main_stage_v_4 & or_tmp_314;
  assign mux_841_nl = MUX_s_1_2_2((and_142_nl), and_tmp_103, or_cse);
  assign nor_573_nl = ~((cfg_precision_1_sva_st_71[1]) | (~ nor_tmp_260));
  assign mux_846_nl = MUX_s_1_2_2((nor_573_nl), nor_tmp_260, cfg_precision_1_sva_st_71[0]);
  assign mux_847_nl = MUX_s_1_2_2((mux_846_nl), main_stage_v_4, and_811_cse);
  assign mux_848_nl = MUX_s_1_2_2((mux_847_nl), mux_845_cse, or_cse);
  assign mux_854_nl = MUX_s_1_2_2(mux_tmp_301, or_tmp_363, or_cse);
  assign or_1113_nl = lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
      | lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
      | (~ and_tmp_108);
  assign mux_855_nl = MUX_s_1_2_2((or_1113_nl), nand_tmp_22, or_cse);
  assign and_1089_nl = or_1857_cse & ((~ FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_2_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_2_sva_7));
  assign mux_1249_nl = MUX_s_1_2_2((and_1089_nl), or_tmp_1720, and_1140_cse);
  assign mux_1250_nl = MUX_s_1_2_2((mux_1249_nl), or_tmp_1720, IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp);
  assign and_147_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 & or_1857_cse & lut_lookup_else_1_slc_32_mdf_2_sva_7
      & main_stage_v_3;
  assign mux_859_nl = MUX_s_1_2_2(and_tmp_108, (and_147_nl), or_cse);
  assign mux_861_nl = MUX_s_1_2_2(mux_805_cse, and_tmp_6, or_cse);
  assign mux_870_nl = MUX_s_1_2_2(nor_564_cse, main_stage_v_3, or_1857_cse);
  assign and_1158_nl = (mux_870_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign mux_875_nl = MUX_s_1_2_2(or_tmp_993, (~ mux_755_cse), lut_lookup_3_if_else_slc_32_svs_8);
  assign or_1142_nl = (~ lut_lookup_3_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3
      | lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign mux_876_nl = MUX_s_1_2_2((mux_875_nl), or_tmp_993, or_1142_nl);
  assign mux_877_nl = MUX_s_1_2_2((mux_876_nl), or_978_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_878_nl = MUX_s_1_2_2((~ (mux_877_nl)), (and_1158_nl), or_cse);
  assign and_149_nl = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & lut_lookup_3_if_else_slc_32_svs_7
      & mux_tmp_704;
  assign mux_880_nl = MUX_s_1_2_2((and_149_nl), main_stage_v_3, or_1857_cse);
  assign and_1156_nl = (mux_880_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign and_808_nl = lut_lookup_3_if_else_slc_32_svs_st_5 & lut_lookup_3_if_else_slc_32_svs_8;
  assign mux_885_nl = MUX_s_1_2_2((~ or_tmp_993), mux_755_cse, and_808_nl);
  assign mux_886_nl = MUX_s_1_2_2((mux_885_nl), nor_612_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_887_nl = MUX_s_1_2_2((mux_886_nl), (and_1156_nl), or_cse);
  assign nor_551_nl = ~((~ lut_lookup_3_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | (~ lut_lookup_3_if_else_else_else_if_acc_itm_3_1) | (~ lut_lookup_3_if_else_slc_32_svs_7)
      | lut_lookup_if_else_else_slc_10_mdf_3_sva_3 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | (~ and_tmp_14));
  assign nor_552_nl = ~((~ lut_lookup_else_else_else_asn_mdf_3_sva_st_3) | cfg_lut_le_function_1_sva_st_42
      | (~ lut_lookup_if_else_else_else_asn_mdf_3_sva_2) | lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3
      | lut_lookup_if_else_else_slc_10_mdf_3_sva_4 | (~(lut_lookup_3_if_else_slc_32_svs_8
      & IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 & lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2
      & lut_lookup_3_if_else_slc_32_svs_st_5 & main_stage_v_4 & or_tmp_314)));
  assign mux_895_nl = MUX_s_1_2_2((nor_552_nl), (nor_551_nl), or_cse);
  assign and_152_nl = lut_lookup_else_else_else_asn_mdf_3_sva_4 & lut_lookup_else_else_else_asn_mdf_3_sva_st_3
      & lut_lookup_else_else_slc_32_mdf_3_sva_8 & cfg_lut_le_function_1_sva_st_42
      & IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 & main_stage_v_4 & or_tmp_314;
  assign mux_896_nl = MUX_s_1_2_2((and_152_nl), and_tmp_113, or_cse);
  assign nor_549_nl = ~((cfg_precision_1_sva_st_71[1]) | (~ nor_tmp_281));
  assign mux_901_nl = MUX_s_1_2_2((nor_549_nl), nor_tmp_281, cfg_precision_1_sva_st_71[0]);
  assign mux_902_nl = MUX_s_1_2_2((mux_901_nl), main_stage_v_4, and_811_cse);
  assign mux_903_nl = MUX_s_1_2_2((mux_902_nl), mux_900_cse, or_cse);
  assign mux_910_nl = MUX_s_1_2_2(or_tmp_573, or_tmp_395, or_cse);
  assign or_1183_nl = lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
      | lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
      | (~ and_tmp_119);
  assign mux_912_nl = MUX_s_1_2_2((or_1183_nl), or_tmp_1181, or_cse);
  assign nor_827_nl = ~(nor_792_cse | (~ FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_3_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_3_sva_7));
  assign nand_102_nl = ~(or_1857_cse & ((~ FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5) |
      FpMantRNE_49U_24U_2_else_carry_3_sva_2 | (~ lut_lookup_else_1_slc_32_mdf_3_sva_7)));
  assign or_2025_nl = and_1139_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp;
  assign mux_1251_nl = MUX_s_1_2_2((nand_102_nl), (nor_827_nl), or_2025_nl);
  assign and_158_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 & lut_lookup_else_1_slc_32_mdf_3_sva_7
      & and_tmp_6;
  assign mux_916_nl = MUX_s_1_2_2(and_tmp_119, (and_158_nl), or_cse);
  assign nor_544_nl = ~((cfg_precision_1_sva_st_71[0]) | (~((cfg_precision_1_sva_st_71[1])
      & main_stage_v_4)));
  assign mux_1284_nl = MUX_s_1_2_2(main_stage_v_4, (nor_544_nl), or_1202_cse);
  assign and_1176_nl = (mux_1284_nl) & (~ cfg_lut_le_function_1_sva_st_42);
  assign mux_926_nl = MUX_s_1_2_2((and_1176_nl), (~ mux_745_cse), or_cse);
  assign nor_540_nl = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (~ FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6)
      | lut_lookup_if_else_else_slc_10_mdf_sva_3 | (~(lut_lookup_4_if_else_slc_32_svs_7
      & mux_tmp_704)));
  assign mux_1271_nl = MUX_s_1_2_2((nor_540_nl), main_stage_v_3, or_1857_cse);
  assign and_1153_nl = (mux_1271_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign mux_933_nl = MUX_s_1_2_2(or_tmp_993, (~ mux_755_cse), lut_lookup_4_if_else_slc_32_svs_8);
  assign or_1213_nl = (~ lut_lookup_4_if_else_slc_32_svs_st_5) | lut_lookup_if_else_else_slc_10_mdf_sva_st_3
      | lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign mux_934_nl = MUX_s_1_2_2((mux_933_nl), or_tmp_993, or_1213_nl);
  assign mux_935_nl = MUX_s_1_2_2((mux_934_nl), or_978_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_936_nl = MUX_s_1_2_2((~ (mux_935_nl)), (and_1153_nl), or_cse);
  assign and_160_nl = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & lut_lookup_4_if_else_slc_32_svs_7
      & mux_tmp_704;
  assign mux_1270_nl = MUX_s_1_2_2((and_160_nl), main_stage_v_3, or_1857_cse);
  assign and_1151_nl = (mux_1270_nl) & (~ cfg_lut_le_function_1_sva_st_41);
  assign and_804_nl = lut_lookup_4_if_else_slc_32_svs_st_5 & lut_lookup_4_if_else_slc_32_svs_8;
  assign mux_943_nl = MUX_s_1_2_2((~ or_tmp_993), mux_755_cse, and_804_nl);
  assign mux_944_nl = MUX_s_1_2_2((mux_943_nl), nor_612_cse, cfg_lut_le_function_1_sva_st_42);
  assign mux_945_nl = MUX_s_1_2_2((mux_944_nl), (and_1151_nl), or_cse);
  assign or_2087_nl = (cfg_precision_1_sva_8!=2'b10) | (cfg_precision_1_sva_st_71[0]);
  assign mux_1283_nl = MUX_s_1_2_2(nor_526_cse, main_stage_v_4, or_2087_nl);
  assign and_1174_nl = (mux_1283_nl) & (~ cfg_lut_le_function_1_sva_st_42);
  assign mux_953_nl = MUX_s_1_2_2((and_1174_nl), mux_771_cse, or_cse);
  assign nor_528_nl = ~((~ lut_lookup_4_if_else_else_else_else_acc_itm_32_1) | cfg_lut_le_function_1_sva_st_41
      | (~ lut_lookup_4_if_else_else_else_if_acc_itm_3_1) | (~ lut_lookup_4_if_else_slc_32_svs_7)
      | lut_lookup_if_else_else_slc_10_mdf_sva_3 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | (~ and_tmp_19));
  assign nor_529_nl = ~(cfg_lut_le_function_1_sva_st_42 | (~ lut_lookup_if_else_else_else_asn_mdf_sva_2)
      | (~ IsNaN_8U_23U_6_land_lpi_1_dfm_6) | (~ lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2)
      | (~ lut_lookup_else_else_else_asn_mdf_sva_st_3) | lut_lookup_if_else_else_slc_10_mdf_sva_4
      | lut_lookup_if_else_else_slc_10_mdf_sva_st_3 | (~(lut_lookup_4_if_else_slc_32_svs_8
      & lut_lookup_4_if_else_slc_32_svs_st_5 & main_stage_v_4 & or_tmp_314)));
  assign mux_954_nl = MUX_s_1_2_2((nor_529_nl), (nor_528_nl), or_cse);
  assign and_163_nl = lut_lookup_else_else_else_asn_mdf_sva_4 & lut_lookup_else_else_slc_32_mdf_sva_8
      & cfg_lut_le_function_1_sva_st_42 & IsNaN_8U_23U_6_land_lpi_1_dfm_6 & lut_lookup_else_else_else_asn_mdf_sva_st_3
      & main_stage_v_4 & or_tmp_314;
  assign mux_955_nl = MUX_s_1_2_2((and_163_nl), and_tmp_124, or_cse);
  assign mux_949_nl = MUX_s_1_2_2(nor_526_cse, main_stage_v_4, cfg_precision_1_sva_st_71[0]);
  assign and_166_nl = cfg_lut_le_function_1_sva_st_42 & IsNaN_8U_23U_6_land_lpi_1_dfm_6
      & lut_lookup_else_else_slc_32_mdf_sva_8 & (mux_949_nl);
  assign mux_961_nl = MUX_s_1_2_2((and_166_nl), main_stage_v_4, and_811_cse);
  assign mux_962_nl = MUX_s_1_2_2((mux_961_nl), mux_959_cse, or_cse);
  assign mux_969_nl = MUX_s_1_2_2(or_tmp_623, or_tmp_427, or_cse);
  assign or_1252_nl = lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3
      | lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3
      | (~ and_tmp_131);
  assign mux_971_nl = MUX_s_1_2_2((or_1252_nl), or_tmp_1250, or_cse);
  assign nor_825_nl = ~(nor_792_cse | (~ FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_sva_7));
  assign nand_nl = ~(or_1857_cse & ((~ FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5) | FpMantRNE_49U_24U_2_else_carry_sva_2
      | (~ lut_lookup_else_1_slc_32_mdf_sva_7)));
  assign or_2035_nl = and_1138_cse | IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp;
  assign mux_1252_nl = MUX_s_1_2_2((nand_nl), (nor_825_nl), or_2035_nl);
  assign mux_975_nl = MUX_s_1_2_2(and_tmp_131, and_tmp_130, or_cse);
  assign nor_518_nl = ~((~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_1_if_else_else_acc_itm_10 | (~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7
      & lut_lookup_1_if_else_slc_32_svs_6 & or_66_cse)));
  assign nor_519_nl = ~(nor_792_cse | (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_1_sva_3
      | (~ lut_lookup_1_if_else_slc_32_svs_7));
  assign nor_521_nl = ~((~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_1_sva_3
      | (~ lut_lookup_1_if_else_slc_32_svs_7));
  assign nor_315_nl = ~(cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6));
  assign mux_980_nl = MUX_s_1_2_2((nor_521_nl), (nor_519_nl), nor_315_nl);
  assign mux_981_nl = MUX_s_1_2_2((mux_980_nl), (nor_518_nl), or_cse);
  assign mux_986_nl = MUX_s_1_2_2(mux_851_cse, and_178_cse, or_cse);
  assign and_179_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & lut_lookup_1_if_else_slc_32_svs_6
      & mux_tmp_655;
  assign mux_1266_nl = MUX_s_1_2_2((and_179_nl), main_stage_v_2, or_66_cse);
  assign and_1147_nl = (mux_1266_nl) & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_995_nl = MUX_s_1_2_2(mux_789_cse, (and_1147_nl), or_cse);
  assign nor_512_nl = ~((~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_2_if_else_else_acc_itm_10 | (~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      & lut_lookup_2_if_else_slc_32_svs_6 & or_66_cse)));
  assign nor_513_nl = ~(nor_792_cse | (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_2_sva_3
      | (~ lut_lookup_2_if_else_slc_32_svs_7));
  assign nor_515_nl = ~((~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_2_sva_3
      | (~ lut_lookup_2_if_else_slc_32_svs_7));
  assign nor_324_nl = ~(cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6));
  assign mux_996_nl = MUX_s_1_2_2((nor_515_nl), (nor_513_nl), nor_324_nl);
  assign mux_997_nl = MUX_s_1_2_2((mux_996_nl), (nor_512_nl), or_cse);
  assign and_193_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & lut_lookup_2_if_else_slc_32_svs_6
      & mux_tmp_655;
  assign mux_1268_nl = MUX_s_1_2_2((and_193_nl), main_stage_v_2, or_66_cse);
  assign and_1149_nl = (mux_1268_nl) & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_1013_nl = MUX_s_1_2_2(mux_845_cse, (and_1149_nl), or_cse);
  assign nor_506_nl = ~((~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_3_if_else_else_acc_itm_10 | (~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      & lut_lookup_3_if_else_slc_32_svs_6 & or_66_cse)));
  assign nor_507_nl = ~(nor_792_cse | (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_3_sva_3
      | (~ lut_lookup_3_if_else_slc_32_svs_7));
  assign nor_509_nl = ~((~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_3_sva_3
      | (~ lut_lookup_3_if_else_slc_32_svs_7));
  assign nor_334_nl = ~(cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6));
  assign mux_1014_nl = MUX_s_1_2_2((nor_509_nl), (nor_507_nl), nor_334_nl);
  assign mux_1015_nl = MUX_s_1_2_2((mux_1014_nl), (nor_506_nl), or_cse);
  assign and_204_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & lut_lookup_3_if_else_slc_32_svs_6
      & mux_tmp_655;
  assign mux_1267_nl = MUX_s_1_2_2((and_204_nl), main_stage_v_2, or_66_cse);
  assign and_1148_nl = (mux_1267_nl) & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_1031_nl = MUX_s_1_2_2(mux_900_cse, (and_1148_nl), or_cse);
  assign nor_500_nl = ~((~ main_stage_v_2) | reg_cfg_lut_le_function_1_sva_st_20_cse
      | lut_lookup_4_if_else_else_acc_itm_10 | (~(IsNaN_8U_23U_1_land_lpi_1_dfm_7
      & lut_lookup_4_if_else_slc_32_svs_6 & or_66_cse)));
  assign nor_501_nl = ~(nor_792_cse | (~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_sva_3
      | (~ lut_lookup_4_if_else_slc_32_svs_7));
  assign nor_503_nl = ~((~ main_stage_v_3) | lut_lookup_if_else_else_slc_10_mdf_sva_3
      | (~ lut_lookup_4_if_else_slc_32_svs_7));
  assign nor_342_nl = ~(cfg_lut_le_function_1_sva_st_41 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | (~ FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6));
  assign mux_1032_nl = MUX_s_1_2_2((nor_503_nl), (nor_501_nl), nor_342_nl);
  assign mux_1033_nl = MUX_s_1_2_2((mux_1032_nl), (nor_500_nl), or_cse);
  assign and_215_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & lut_lookup_4_if_else_slc_32_svs_6
      & mux_tmp_655;
  assign mux_nl = MUX_s_1_2_2((and_215_nl), main_stage_v_2, or_66_cse);
  assign and_1146_nl = (mux_nl) & reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign mux_1049_nl = MUX_s_1_2_2(mux_959_cse, (and_1146_nl), or_cse);
  assign mux_1051_nl = MUX_s_1_2_2(and_tmp_6, mux_982_cse, or_cse);
  assign mux_1055_nl = MUX_s_1_2_2(mux_793_cse, and_42_cse, or_cse);
  assign nor_495_nl = ~(and_794_cse | and_795_cse | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_lut_in_rsci_bawt));
  assign nor_496_nl = ~((~ reg_cfg_lut_le_function_1_sva_st_19_cse) | (~ main_stage_v_1)
      | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6);
  assign nor_497_nl = ~((~(IsNaN_8U_23U_4_nor_itm_2 | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2
      | (~ reg_cfg_lut_le_function_1_sva_st_19_cse))) | (~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6);
  assign mux_1057_nl = MUX_s_1_2_2((nor_497_nl), (nor_496_nl), IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4);
  assign mux_1058_nl = MUX_s_1_2_2((mux_1057_nl), (nor_495_nl), or_cse);
  assign nor_493_nl = ~(and_795_cse | (cfg_precision_rsci_d!=2'b10) | (~(cfg_lut_le_function_rsci_d
      & chn_lut_in_rsci_bawt)));
  assign nor_494_nl = ~((~ main_stage_v_1) | (~ reg_cfg_lut_le_function_1_sva_st_19_cse)
      | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10) | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4);
  assign mux_1059_nl = MUX_s_1_2_2((nor_494_nl), (nor_493_nl), or_cse);
  assign nor_491_nl = ~(((~ IsNaN_8U_23U_3_nor_8_tmp) & (chn_lut_in_rsci_d_mxwt[30:23]==8'b11111111)
      & cfg_lut_le_function_rsci_d) | (cfg_precision_rsci_d!=2'b10) | (~ chn_lut_in_rsci_bawt));
  assign nor_492_nl = ~((reg_cfg_lut_le_function_1_sva_st_19_cse & IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4)
      | (~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign mux_1060_nl = MUX_s_1_2_2((nor_492_nl), (nor_491_nl), or_cse);
  assign nor_489_nl = ~(and_789_cse | and_795_cse | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_lut_in_rsci_bawt));
  assign nor_490_nl = ~((~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_5);
  assign mux_1061_nl = MUX_s_1_2_2((nor_490_nl), (nor_489_nl), or_cse);
  assign nor_487_nl = ~(and_787_cse | or_tmp_1360);
  assign nor_488_nl = ~((reg_cfg_precision_1_sva_st_12_cse_1!=2'b10) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 | (~ main_stage_v_1));
  assign mux_1062_nl = MUX_s_1_2_2((nor_488_nl), (nor_487_nl), or_cse);
  assign nor_485_nl = ~(and_789_cse | and_787_cse | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_lut_in_rsci_bawt));
  assign nor_486_nl = ~((~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 | IsNaN_8U_23U_8_land_2_lpi_1_dfm_5);
  assign mux_1063_nl = MUX_s_1_2_2((nor_486_nl), (nor_485_nl), or_cse);
  assign nor_483_nl = ~(and_784_cse | or_tmp_1360);
  assign nor_484_nl = ~((~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4);
  assign mux_1064_nl = MUX_s_1_2_2((nor_484_nl), (nor_483_nl), or_cse);
  assign nor_480_nl = ~(and_789_cse | and_784_cse | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_lut_in_rsci_bawt));
  assign nor_481_nl = ~((~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 | nor_482_cse);
  assign mux_1066_nl = MUX_s_1_2_2((nor_481_nl), (nor_480_nl), or_cse);
  assign nor_475_nl = ~(and_794_cse | and_780_cse | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_lut_in_rsci_bawt));
  assign nor_476_nl = ~((~ reg_cfg_lut_le_function_1_sva_st_19_cse) | (~ main_stage_v_1)
      | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10) | IsNaN_8U_23U_1_land_lpi_1_dfm_6);
  assign nor_477_nl = ~((~(IsNaN_8U_23U_4_nor_3_itm_2 | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2
      | (~ reg_cfg_lut_le_function_1_sva_st_19_cse))) | (~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | IsNaN_8U_23U_1_land_lpi_1_dfm_6);
  assign mux_1068_nl = MUX_s_1_2_2((nor_477_nl), (nor_476_nl), reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse);
  assign mux_1069_nl = MUX_s_1_2_2((mux_1068_nl), (nor_475_nl), or_cse);
  assign nor_472_nl = ~((~(cfg_lut_le_function_rsci_d & chn_lut_in_rsci_bawt & (cfg_precision_rsci_d==2'b10)))
      | IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0);
  assign nor_473_nl = ~(reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse | (~ main_stage_v_1)
      | (~ reg_cfg_lut_le_function_1_sva_st_19_cse) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign mux_1070_nl = MUX_s_1_2_2((nor_473_nl), (nor_472_nl), or_cse);
  assign nor_470_nl = ~(((~ IsNaN_8U_23U_3_nor_6_tmp) & (chn_lut_in_rsci_d_mxwt[126:119]==8'b11111111)
      & cfg_lut_le_function_rsci_d) | (cfg_precision_rsci_d!=2'b10) | (~ chn_lut_in_rsci_bawt));
  assign nor_471_nl = ~((reg_cfg_lut_le_function_1_sva_st_19_cse & reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse)
      | (~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10));
  assign mux_1071_nl = MUX_s_1_2_2((nor_471_nl), (nor_470_nl), or_cse);
  assign nor_467_nl = ~(and_789_cse | and_780_cse | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_lut_in_rsci_bawt));
  assign nor_468_nl = ~((~ main_stage_v_1) | (reg_cfg_precision_1_sva_st_12_cse_1!=2'b10)
      | reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse | nor_469_cse);
  assign mux_1073_nl = MUX_s_1_2_2((nor_468_nl), (nor_467_nl), or_cse);
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_1_nl = MUX_v_6_2_2(6'b000000,
      (IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva[5:0]), lut_lookup_1_else_else_else_if_acc_itm_3_1);
  assign and_219_nl = lut_lookup_1_if_else_slc_32_svs_6 & main_stage_v_2 & or_66_cse;
  assign nor_463_nl = ~((~ lut_lookup_1_if_else_slc_32_svs_6) | lut_lookup_1_if_else_else_acc_itm_10
      | (~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & main_stage_v_2 & or_66_cse)));
  assign mux_1075_nl = MUX_s_1_2_2((nor_463_nl), (and_219_nl), reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign and_220_nl = lut_lookup_else_else_slc_32_mdf_1_sva_7 & main_stage_v_3 &
      or_1857_cse;
  assign nor_464_nl = ~((~ lut_lookup_1_if_else_slc_32_svs_7) | lut_lookup_if_else_else_slc_10_mdf_1_sva_3
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (~ and_tmp_5));
  assign mux_1076_nl = MUX_s_1_2_2((nor_464_nl), (and_220_nl), cfg_lut_le_function_1_sva_st_41);
  assign mux_1077_nl = MUX_s_1_2_2((mux_1076_nl), (mux_1075_nl), or_cse);
  assign and_221_nl = lut_lookup_1_else_else_else_if_acc_itm_3_1 & reg_cfg_lut_le_function_1_sva_st_20_cse
      & lut_lookup_1_if_else_slc_32_svs_6 & IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & main_stage_v_2
      & or_66_cse;
  assign mux_1078_nl = MUX_s_1_2_2(and_tmp_92, (and_221_nl), or_cse);
  assign or_1431_nl = (~ lut_lookup_else_1_slc_32_mdf_1_sva_6) | (lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])
      | (~ and_tmp_61);
  assign mux_1079_nl = MUX_s_1_2_2(or_tmp_1043, (or_1431_nl), or_cse);
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_3_nl = MUX_v_6_2_2(6'b000000,
      (IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva[5:0]), lut_lookup_2_else_else_else_if_acc_itm_3_1);
  assign and_222_nl = lut_lookup_2_if_else_slc_32_svs_6 & mux_tmp_655;
  assign nor_459_nl = ~(lut_lookup_2_if_else_else_acc_itm_10 | (~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      & lut_lookup_2_if_else_slc_32_svs_6 & mux_tmp_655)));
  assign mux_1081_nl = MUX_s_1_2_2((nor_459_nl), (and_222_nl), reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign and_224_nl = lut_lookup_else_else_slc_32_mdf_2_sva_7 & mux_tmp_704;
  assign mux_1083_nl = MUX_s_1_2_2(nor_588_cse, (and_224_nl), cfg_lut_le_function_1_sva_st_41);
  assign mux_1084_nl = MUX_s_1_2_2((mux_1083_nl), (mux_1081_nl), or_cse);
  assign and_226_nl = lut_lookup_2_if_else_slc_32_svs_6 & IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      & lut_lookup_2_else_else_else_if_acc_itm_3_1 & reg_cfg_lut_le_function_1_sva_st_20_cse
      & main_stage_v_2 & or_66_cse;
  assign mux_1085_nl = MUX_s_1_2_2(and_tmp_103, (and_226_nl), or_cse);
  assign or_1440_nl = (lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])
      | (~(lut_lookup_else_1_slc_32_mdf_2_sva_6 & IsNaN_8U_23U_7_land_2_lpi_1_dfm_6
      & mux_tmp_655));
  assign mux_1086_nl = MUX_s_1_2_2(nand_tmp_22, (or_1440_nl), or_cse);
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_5_nl = MUX_v_6_2_2(6'b000000,
      (IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva[5:0]), lut_lookup_3_else_else_else_if_acc_itm_3_1);
  assign and_228_nl = lut_lookup_3_if_else_slc_32_svs_6 & mux_tmp_655;
  assign nor_455_nl = ~(lut_lookup_3_if_else_else_acc_itm_10 | (~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      & lut_lookup_3_if_else_slc_32_svs_6 & mux_tmp_655)));
  assign mux_1088_nl = MUX_s_1_2_2((nor_455_nl), (and_228_nl), reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign and_230_nl = lut_lookup_else_else_slc_32_mdf_3_sva_7 & mux_tmp_704;
  assign mux_1090_nl = MUX_s_1_2_2(nor_564_cse, (and_230_nl), cfg_lut_le_function_1_sva_st_41);
  assign mux_1091_nl = MUX_s_1_2_2((mux_1090_nl), (mux_1088_nl), or_cse);
  assign and_232_nl = lut_lookup_3_if_else_slc_32_svs_6 & IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      & lut_lookup_3_else_else_else_if_acc_itm_3_1 & reg_cfg_lut_le_function_1_sva_st_20_cse
      & main_stage_v_2 & or_66_cse;
  assign mux_1092_nl = MUX_s_1_2_2(and_tmp_113, (and_232_nl), or_cse);
  assign or_1450_nl = (~ lut_lookup_else_1_slc_32_mdf_3_sva_6) | (lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])
      | (~ and_tmp_69);
  assign mux_1093_nl = MUX_s_1_2_2(or_tmp_1181, (or_1450_nl), or_cse);
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_7_nl = MUX_v_6_2_2(6'b000000,
      (IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva[5:0]), lut_lookup_4_else_else_else_if_acc_itm_3_1);
  assign and_233_nl = lut_lookup_4_if_else_slc_32_svs_6 & main_stage_v_2 & or_66_cse;
  assign nor_453_nl = ~((~ lut_lookup_4_if_else_slc_32_svs_6) | lut_lookup_4_if_else_else_acc_itm_10
      | (~(IsNaN_8U_23U_1_land_lpi_1_dfm_7 & main_stage_v_2 & or_66_cse)));
  assign mux_1094_nl = MUX_s_1_2_2((nor_453_nl), (and_233_nl), reg_cfg_lut_le_function_1_sva_st_20_cse);
  assign and_235_nl = lut_lookup_else_else_slc_32_mdf_sva_7 & main_stage_v_3 & or_1857_cse;
  assign nor_454_nl = ~((~ lut_lookup_4_if_else_slc_32_svs_7) | lut_lookup_if_else_else_slc_10_mdf_sva_3
      | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (~ and_tmp_19));
  assign mux_1095_nl = MUX_s_1_2_2((nor_454_nl), (and_235_nl), cfg_lut_le_function_1_sva_st_41);
  assign mux_1096_nl = MUX_s_1_2_2((mux_1095_nl), (mux_1094_nl), or_cse);
  assign and_236_nl = reg_cfg_lut_le_function_1_sva_st_20_cse & IsNaN_8U_23U_1_land_lpi_1_dfm_7
      & lut_lookup_4_else_else_else_if_acc_itm_3_1 & lut_lookup_4_if_else_slc_32_svs_6
      & main_stage_v_2 & or_66_cse;
  assign mux_1097_nl = MUX_s_1_2_2(and_tmp_124, (and_236_nl), or_cse);
  assign or_1458_nl = (lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8])
      | (~(lut_lookup_else_1_slc_32_mdf_sva_6 & IsNaN_8U_23U_7_land_lpi_1_dfm_6 &
      main_stage_v_2 & or_66_cse));
  assign mux_1098_nl = MUX_s_1_2_2(or_tmp_1250, (or_1458_nl), or_cse);
  assign nand_33_nl = ~(main_stage_v_1 & lut_lookup_1_if_else_slc_32_svs_5);
  assign or_1830_nl = reg_cfg_lut_le_function_1_sva_st_20_cse | not_tmp_800;
  assign mux_1099_nl = MUX_s_1_2_2((or_1830_nl), (nand_33_nl), or_cse);
  assign mux_1100_nl = MUX_s_1_2_2(or_tmp_1450, (mux_1099_nl), FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign or_1460_nl = nor_190_cse | reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign mux_1101_nl = MUX_s_1_2_2((mux_1100_nl), or_tmp_1450, or_1460_nl);
  assign mux_1103_nl = MUX_s_1_2_2(and_42_cse, mux_tmp_1101, or_cse);
  assign nor_451_nl = ~(reg_cfg_lut_le_function_1_sva_st_19_cse | (~(FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5
      & or_26_cse & main_stage_v_1 & lut_lookup_2_if_else_slc_32_svs_5)));
  assign and_774_nl = lut_lookup_2_if_else_slc_32_svs_6 & IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      & (~ reg_cfg_lut_le_function_1_sva_st_20_cse) & and_42_cse;
  assign mux_1104_nl = MUX_s_1_2_2((and_774_nl), (nor_451_nl), or_cse);
  assign nor_450_nl = ~((~ main_stage_v_1) | (~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5)
      | reg_cfg_lut_le_function_1_sva_st_19_cse | (~(or_26_cse & lut_lookup_3_if_else_slc_32_svs_5)));
  assign and_773_nl = lut_lookup_3_if_else_slc_32_svs_6 & IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      & (~ reg_cfg_lut_le_function_1_sva_st_20_cse) & and_42_cse;
  assign mux_1107_nl = MUX_s_1_2_2((and_773_nl), (nor_450_nl), or_cse);
  assign nor_448_nl = ~((~ main_stage_v_1) | (~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5)
      | reg_cfg_lut_le_function_1_sva_st_19_cse | (~(or_26_cse & lut_lookup_4_if_else_slc_32_svs_5)));
  assign nor_449_nl = ~(reg_cfg_lut_le_function_1_sva_st_20_cse | (~(lut_lookup_4_if_else_slc_32_svs_6
      & IsNaN_8U_23U_1_land_lpi_1_dfm_7 & main_stage_v_2 & or_66_cse)));
  assign mux_1110_nl = MUX_s_1_2_2((nor_449_nl), (nor_448_nl), or_cse);
  assign mux_1112_nl = MUX_s_1_2_2(mux_982_cse, mux_tmp_1104, or_cse);
  assign mux_1118_nl = MUX_s_1_2_2(mux_tmp_1101, and_tmp_178, or_cse);
  assign nl_z_out_4 = conv_u2u_8_9(FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp) + 9'b110000001;
  assign z_out_4 = nl_z_out_4[8:0];
  assign nl_z_out_5 = conv_u2u_8_9(FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7) + 9'b110000001;
  assign z_out_5 = nl_z_out_5[8:0];
  assign nl_z_out_6 = conv_u2u_8_9(FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7) + 9'b110000001;
  assign z_out_6 = nl_z_out_6[8:0];
  assign nl_z_out_7 = conv_u2u_8_9(FpAdd_8U_23U_o_expo_lpi_1_dfm_7) + 9'b110000001;
  assign z_out_7 = nl_z_out_7[8:0];
  assign nand_113_nl = ~(lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 &
      mux_tmp_1247);
  assign or_2088_nl = lut_lookup_else_if_lor_5_lpi_1_dfm_6 | lut_lookup_1_else_if_else_if_acc_itm_3_1
      | (~ mux_tmp_1247);
  assign mux_1289_nl = MUX_s_1_2_2((or_2088_nl), (nand_113_nl), lut_lookup_unequal_tmp_13);
  assign nand_114_nl = ~(lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 &
      mux_tmp_1247);
  assign mux_1288_nl = MUX_s_1_2_2((nand_114_nl), (mux_1289_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_else_2_else_else_else_and_4_nl = (fsm_output[1]) & (mux_1288_nl);
  assign lut_lookup_else_2_if_mux_31_nl = MUX_s_1_2_2(cfg_lut_oflow_priority_1_sva_10,
      lut_lookup_le_miss_1_sva, lut_lookup_else_2_else_else_else_and_4_nl);
  assign z_out = MUX_s_1_2_2(lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0, (lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[0]),
      lut_lookup_else_2_if_mux_31_nl);
  assign nand_115_nl = ~(lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 &
      mux_tmp_1250);
  assign or_2089_nl = lut_lookup_else_if_lor_6_lpi_1_dfm_6 | lut_lookup_2_else_if_else_if_acc_itm_3_1
      | (~ mux_tmp_1250);
  assign mux_1292_nl = MUX_s_1_2_2((or_2089_nl), (nand_115_nl), lut_lookup_else_unequal_tmp_13);
  assign nand_116_nl = ~(lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 &
      mux_tmp_1250);
  assign mux_1291_nl = MUX_s_1_2_2((nand_116_nl), (mux_1292_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_else_2_else_else_else_and_5_nl = (fsm_output[1]) & (mux_1291_nl);
  assign lut_lookup_else_2_if_mux_32_nl = MUX_s_1_2_2(cfg_lut_oflow_priority_1_sva_10,
      lut_lookup_le_miss_2_sva, lut_lookup_else_2_else_else_else_and_5_nl);
  assign z_out_1 = MUX_s_1_2_2(lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0, (lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[0]),
      lut_lookup_else_2_if_mux_32_nl);
  assign nand_117_nl = ~(lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 &
      mux_tmp_1253);
  assign or_2090_nl = lut_lookup_else_if_lor_7_lpi_1_dfm_6 | lut_lookup_3_else_if_else_if_acc_itm_3_1
      | (~ mux_tmp_1253);
  assign mux_1295_nl = MUX_s_1_2_2((or_2090_nl), (nand_117_nl), lut_lookup_else_unequal_tmp_13);
  assign nand_118_nl = ~(lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 &
      mux_tmp_1253);
  assign mux_1294_nl = MUX_s_1_2_2((nand_118_nl), (mux_1295_nl), cfg_lut_le_function_1_sva_10);
  assign lut_lookup_else_2_else_else_else_and_6_nl = (fsm_output[1]) & (mux_1294_nl);
  assign lut_lookup_else_2_if_mux_33_nl = MUX_s_1_2_2(cfg_lut_oflow_priority_1_sva_10,
      lut_lookup_le_miss_3_sva, lut_lookup_else_2_else_else_else_and_6_nl);
  assign z_out_2 = MUX_s_1_2_2(lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0, (lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[0]),
      lut_lookup_else_2_if_mux_33_nl);
  assign nor_882_nl = ~(lut_lookup_else_if_lor_1_lpi_1_dfm_6 | lut_lookup_4_else_if_else_if_acc_itm_3_1
      | (~ mux_tmp_1257));
  assign mux_1298_nl = MUX_s_1_2_2(and_tmp_201, (nor_882_nl), cfg_lut_le_function_1_sva_10);
  assign mux_1297_nl = MUX_s_1_2_2((mux_1298_nl), and_tmp_201, lut_lookup_else_unequal_tmp_13);
  assign lut_lookup_else_2_else_else_else_and_7_nl = (fsm_output[1]) & (~ (mux_1297_nl));
  assign lut_lookup_else_2_if_mux_34_nl = MUX_s_1_2_2(cfg_lut_oflow_priority_1_sva_10,
      lut_lookup_le_miss_sva, lut_lookup_else_2_else_else_else_and_7_nl);
  assign z_out_3 = MUX_s_1_2_2(lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0, (lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[0]),
      lut_lookup_else_2_if_mux_34_nl);

  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function [11:0] MUX1HOT_v_12_5_2;
    input [11:0] input_4;
    input [11:0] input_3;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [4:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | ( input_1 & {12{sel[1]}});
    result = result | ( input_2 & {12{sel[2]}});
    result = result | ( input_3 & {12{sel[3]}});
    result = result | ( input_4 & {12{sel[4]}});
    MUX1HOT_v_12_5_2 = result;
  end
  endfunction


  function [22:0] MUX1HOT_v_23_6_2;
    input [22:0] input_5;
    input [22:0] input_4;
    input [22:0] input_3;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [5:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    result = result | ( input_3 & {23{sel[3]}});
    result = result | ( input_4 & {23{sel[4]}});
    result = result | ( input_5 & {23{sel[5]}});
    MUX1HOT_v_23_6_2 = result;
  end
  endfunction


  function [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function [49:0] MUX1HOT_v_50_4_2;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [3:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | ( input_1 & {50{sel[1]}});
    result = result | ( input_2 & {50{sel[2]}});
    result = result | ( input_3 & {50{sel[3]}});
    MUX1HOT_v_50_4_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    result = result | ( input_4 & {6{sel[4]}});
    result = result | ( input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_5_2;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [4:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    MUX1HOT_v_8_5_2 = result;
  end
  endfunction


  function [8:0] MUX1HOT_v_9_5_2;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [4:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    result = result | ( input_4 & {9{sel[4]}});
    MUX1HOT_v_9_5_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function [34:0] MUX_v_35_2_2;
    input [34:0] input_0;
    input [34:0] input_1;
    input [0:0] sel;
    reg [34:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_35_2_2 = result;
  end
  endfunction


  function [48:0] MUX_v_49_2_2;
    input [48:0] input_0;
    input [48:0] input_1;
    input [0:0] sel;
    reg [48:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_49_2_2 = result;
  end
  endfunction


  function [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_248_1_247;
    input [247:0] vector;
    reg [247:0] tmp;
  begin
    tmp = vector >> 247;
    readslicef_248_1_247 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_24_1_23;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 23;
    readslicef_24_1_23 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function [22:0] signext_23_1;
    input [0:0] vector;
  begin
    signext_23_1= {{22{vector[0]}}, vector};
  end
  endfunction


  function [31:0] signext_32_6;
    input [5:0] vector;
  begin
    signext_32_6= {{26{vector[5]}}, vector};
  end
  endfunction


  function [34:0] signext_35_1;
    input [0:0] vector;
  begin
    signext_35_1= {{34{vector[0]}}, vector};
  end
  endfunction


  function [5:0] signext_6_1;
    input [0:0] vector;
  begin
    signext_6_1= {{5{vector[0]}}, vector};
  end
  endfunction


  function [7:0] signext_8_1;
    input [0:0] vector;
  begin
    signext_8_1= {{7{vector[0]}}, vector};
  end
  endfunction


  function [8:0] signext_9_6;
    input [5:0] vector;
  begin
    signext_9_6= {{3{vector[5]}}, vector};
  end
  endfunction


  function  [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function  [9:0] conv_s2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function  [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function  [6:0] conv_s2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction


  function  [8:0] conv_s2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_9 = {{3{vector[5]}}, vector};
  end
  endfunction


  function  [7:0] conv_s2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_8 = {vector[6], vector};
  end
  endfunction


  function  [8:0] conv_s2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_9 = {vector[7], vector};
  end
  endfunction


  function  [9:0] conv_s2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function  [10:0] conv_s2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_11 = {{3{vector[7]}}, vector};
  end
  endfunction


  function  [9:0] conv_s2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_10 = {vector[8], vector};
  end
  endfunction


  function  [32:0] conv_s2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction


  function  [8:0] conv_u2s_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function  [32:0] conv_u2s_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2s_32_33 =  {1'b0, vector};
  end
  endfunction


  function  [22:0] conv_u2u_1_23 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction


  function  [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function  [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function  [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [23:0] conv_u2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_u2u_23_24 = {1'b0, vector};
  end
  endfunction


  function  [49:0] conv_u2u_49_50 ;
    input [48:0]  vector ;
  begin
    conv_u2u_49_50 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_idx
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_idx (
  nvdla_core_clk, nvdla_core_rstn, chn_lut_in_rsc_z, chn_lut_in_rsc_vz, chn_lut_in_rsc_lz,
      cfg_lut_le_start_rsc_z, cfg_lut_lo_start_rsc_z, cfg_lut_le_index_offset_rsc_z,
      cfg_lut_le_index_select_rsc_z, cfg_lut_lo_index_select_rsc_z, cfg_lut_le_function_rsc_z,
      cfg_lut_uflow_priority_rsc_z, cfg_lut_oflow_priority_rsc_z, cfg_lut_hybrid_priority_rsc_z,
      cfg_precision_rsc_z, chn_lut_out_rsc_z, chn_lut_out_rsc_vz, chn_lut_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_lut_in_rsc_z;
  input chn_lut_in_rsc_vz;
  output chn_lut_in_rsc_lz;
  input [31:0] cfg_lut_le_start_rsc_z;
  input [31:0] cfg_lut_lo_start_rsc_z;
  input [7:0] cfg_lut_le_index_offset_rsc_z;
  input [7:0] cfg_lut_le_index_select_rsc_z;
  input [7:0] cfg_lut_lo_index_select_rsc_z;
  input cfg_lut_le_function_rsc_z;
  input cfg_lut_uflow_priority_rsc_z;
  input cfg_lut_oflow_priority_rsc_z;
  input cfg_lut_hybrid_priority_rsc_z;
  input [1:0] cfg_precision_rsc_z;
  output [323:0] chn_lut_out_rsc_z;
  input chn_lut_out_rsc_vz;
  output chn_lut_out_rsc_lz;


  // Interconnect Declarations
  wire chn_lut_in_rsci_oswt;
  wire chn_lut_in_rsci_oswt_unreg;
  wire chn_lut_out_rsci_oswt;
  wire chn_lut_out_rsci_oswt_unreg;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_IDX_chn_lut_in_rsci_unreg chn_lut_in_rsci_unreg_inst (
      .in_0(chn_lut_in_rsci_oswt_unreg),
      .outsig(chn_lut_in_rsci_oswt)
    );
  SDP_Y_IDX_chn_lut_out_rsci_unreg chn_lut_out_rsci_unreg_inst (
      .in_0(chn_lut_out_rsci_oswt_unreg),
      .outsig(chn_lut_out_rsci_oswt)
    );
  NV_NVDLA_SDP_CORE_Y_idx_core NV_NVDLA_SDP_CORE_Y_idx_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_lut_in_rsc_z(chn_lut_in_rsc_z),
      .chn_lut_in_rsc_vz(chn_lut_in_rsc_vz),
      .chn_lut_in_rsc_lz(chn_lut_in_rsc_lz),
      .cfg_lut_le_start_rsc_z(cfg_lut_le_start_rsc_z),
      .cfg_lut_lo_start_rsc_z(cfg_lut_lo_start_rsc_z),
      .cfg_lut_le_index_offset_rsc_z(cfg_lut_le_index_offset_rsc_z),
      .cfg_lut_le_index_select_rsc_z(cfg_lut_le_index_select_rsc_z),
      .cfg_lut_lo_index_select_rsc_z(cfg_lut_lo_index_select_rsc_z),
      .cfg_lut_le_function_rsc_z(cfg_lut_le_function_rsc_z),
      .cfg_lut_uflow_priority_rsc_z(cfg_lut_uflow_priority_rsc_z),
      .cfg_lut_oflow_priority_rsc_z(cfg_lut_oflow_priority_rsc_z),
      .cfg_lut_hybrid_priority_rsc_z(cfg_lut_hybrid_priority_rsc_z),
      .cfg_precision_rsc_z(cfg_precision_rsc_z),
      .chn_lut_out_rsc_z(chn_lut_out_rsc_z),
      .chn_lut_out_rsc_vz(chn_lut_out_rsc_vz),
      .chn_lut_out_rsc_lz(chn_lut_out_rsc_lz),
      .chn_lut_in_rsci_oswt(chn_lut_in_rsci_oswt),
      .chn_lut_in_rsci_oswt_unreg(chn_lut_in_rsci_oswt_unreg),
      .chn_lut_out_rsci_oswt(chn_lut_out_rsci_oswt),
      .chn_lut_out_rsci_oswt_unreg(chn_lut_out_rsci_oswt_unreg)
    );
endmodule



