// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: HLS_fp32_mul.v

module FP32_MUL_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/FP32_MUL_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module FP32_MUL_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-184
//  Generated date: Fri Jun 16 21:53:54 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    FP32_MUL_chn_o_rsci_unreg
// ------------------------------------------------------------------


module FP32_MUL_chn_o_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP32_MUL_chn_b_rsci_unreg
// ------------------------------------------------------------------


module FP32_MUL_chn_b_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP32_MUL_chn_a_rsci_unreg
// ------------------------------------------------------------------


module FP32_MUL_chn_a_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module HLS_fp32_mul_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for HLS_fp32_mul_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : HLS_fp32_mul_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_staller
// ------------------------------------------------------------------


module HLS_fp32_mul_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_a_rsci_wen_comp, core_wten, chn_b_rsci_wen_comp,
      chn_o_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_a_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_b_rsci_wen_comp;
  input chn_o_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_a_rsci_wen_comp & chn_b_rsci_wen_comp & chn_o_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_dp
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_biwt, chn_o_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_biwt;
  input chn_o_rsci_bdwt;


  // Interconnect Declarations
  reg chn_o_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_bawt = chn_o_rsci_biwt | chn_o_rsci_bcwt;
  assign chn_o_rsci_wen_comp = (~ chn_o_rsci_oswt) | chn_o_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_o_rsci_bcwt <= ~((~(chn_o_rsci_bcwt | chn_o_rsci_biwt)) | chn_o_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, core_wen, core_wten, chn_o_rsci_iswt0,
      chn_o_rsci_ld_core_psct, chn_o_rsci_biwt, chn_o_rsci_bdwt, chn_o_rsci_ld_core_sct,
      chn_o_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  input chn_o_rsci_ld_core_psct;
  output chn_o_rsci_biwt;
  output chn_o_rsci_bdwt;
  output chn_o_rsci_ld_core_sct;
  input chn_o_rsci_vd;


  // Interconnect Declarations
  wire chn_o_rsci_ogwt;
  wire chn_o_rsci_pdswt0;
  reg chn_o_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_pdswt0 = (~ core_wten) & chn_o_rsci_iswt0;
  assign chn_o_rsci_biwt = chn_o_rsci_ogwt & chn_o_rsci_vd;
  assign chn_o_rsci_ogwt = chn_o_rsci_pdswt0 | chn_o_rsci_icwt;
  assign chn_o_rsci_bdwt = chn_o_rsci_oswt & core_wen;
  assign chn_o_rsci_ld_core_sct = chn_o_rsci_ld_core_psct & chn_o_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_icwt <= 1'b0;
    end
    else begin
      chn_o_rsci_icwt <= ~((~(chn_o_rsci_icwt | chn_o_rsci_pdswt0)) | chn_o_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_dp
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsci_oswt, chn_b_rsci_bawt, chn_b_rsci_wen_comp,
      chn_b_rsci_d_mxwt, chn_b_rsci_biwt, chn_b_rsci_bdwt, chn_b_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_b_rsci_oswt;
  output chn_b_rsci_bawt;
  output chn_b_rsci_wen_comp;
  output [31:0] chn_b_rsci_d_mxwt;
  input chn_b_rsci_biwt;
  input chn_b_rsci_bdwt;
  input [31:0] chn_b_rsci_d;


  // Interconnect Declarations
  reg chn_b_rsci_bcwt;
  reg [31:0] chn_b_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_b_rsci_bawt = chn_b_rsci_biwt | chn_b_rsci_bcwt;
  assign chn_b_rsci_wen_comp = (~ chn_b_rsci_oswt) | chn_b_rsci_bawt;
  assign chn_b_rsci_d_mxwt = MUX_v_32_2_2(chn_b_rsci_d, chn_b_rsci_d_bfwt, chn_b_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_b_rsci_bcwt <= 1'b0;
      chn_b_rsci_d_bfwt <= 32'b0;
    end
    else begin
      chn_b_rsci_bcwt <= ~((~(chn_b_rsci_bcwt | chn_b_rsci_biwt)) | chn_b_rsci_bdwt);
      chn_b_rsci_d_bfwt <= chn_b_rsci_d_mxwt;
    end
  end

  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsci_oswt, core_wen, core_wten, chn_b_rsci_iswt0,
      chn_b_rsci_ld_core_psct, chn_b_rsci_biwt, chn_b_rsci_bdwt, chn_b_rsci_ld_core_sct,
      chn_b_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_b_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_b_rsci_iswt0;
  input chn_b_rsci_ld_core_psct;
  output chn_b_rsci_biwt;
  output chn_b_rsci_bdwt;
  output chn_b_rsci_ld_core_sct;
  input chn_b_rsci_vd;


  // Interconnect Declarations
  wire chn_b_rsci_ogwt;
  wire chn_b_rsci_pdswt0;
  reg chn_b_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_b_rsci_pdswt0 = (~ core_wten) & chn_b_rsci_iswt0;
  assign chn_b_rsci_biwt = chn_b_rsci_ogwt & chn_b_rsci_vd;
  assign chn_b_rsci_ogwt = chn_b_rsci_pdswt0 | chn_b_rsci_icwt;
  assign chn_b_rsci_bdwt = chn_b_rsci_oswt & core_wen;
  assign chn_b_rsci_ld_core_sct = chn_b_rsci_ld_core_psct & chn_b_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_b_rsci_icwt <= 1'b0;
    end
    else begin
      chn_b_rsci_icwt <= ~((~(chn_b_rsci_icwt | chn_b_rsci_pdswt0)) | chn_b_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_dp
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, chn_a_rsci_bawt, chn_a_rsci_wen_comp,
      chn_a_rsci_d_mxwt, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  output [31:0] chn_a_rsci_d_mxwt;
  input chn_a_rsci_biwt;
  input chn_a_rsci_bdwt;
  input [31:0] chn_a_rsci_d;


  // Interconnect Declarations
  reg chn_a_rsci_bcwt;
  reg [31:0] chn_a_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_bawt = chn_a_rsci_biwt | chn_a_rsci_bcwt;
  assign chn_a_rsci_wen_comp = (~ chn_a_rsci_oswt) | chn_a_rsci_bawt;
  assign chn_a_rsci_d_mxwt = MUX_v_32_2_2(chn_a_rsci_d, chn_a_rsci_d_bfwt, chn_a_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_bcwt <= 1'b0;
      chn_a_rsci_d_bfwt <= 32'b0;
    end
    else begin
      chn_a_rsci_bcwt <= ~((~(chn_a_rsci_bcwt | chn_a_rsci_biwt)) | chn_a_rsci_bdwt);
      chn_a_rsci_d_bfwt <= chn_a_rsci_d_mxwt;
    end
  end

  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct,
      core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  input chn_a_rsci_ld_core_psct;
  input core_wten;
  output chn_a_rsci_biwt;
  output chn_a_rsci_bdwt;
  output chn_a_rsci_ld_core_sct;
  input chn_a_rsci_vd;


  // Interconnect Declarations
  wire chn_a_rsci_ogwt;
  wire chn_a_rsci_pdswt0;
  reg chn_a_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_pdswt0 = (~ core_wten) & chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & chn_a_rsci_vd;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | chn_a_rsci_icwt;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & chn_a_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_icwt <= 1'b0;
    end
    else begin
      chn_a_rsci_icwt <= ~((~(chn_a_rsci_icwt | chn_a_rsci_pdswt0)) | chn_a_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_o_rsci
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_o_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_o_rsci_oswt,
      core_wen, core_wten, chn_o_rsci_iswt0, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_ld_core_psct, chn_o_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [31:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_ld_core_psct;
  input [31:0] chn_o_rsci_d;


  // Interconnect Declarations
  wire chn_o_rsci_biwt;
  wire chn_o_rsci_bdwt;
  wire chn_o_rsci_ld_core_sct;
  wire chn_o_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  FP32_MUL_mgc_out_stdreg_wait_v1 #(.rscid(32'sd3),
  .width(32'sd32)) chn_o_rsci (
      .ld(chn_o_rsci_ld_core_sct),
      .vd(chn_o_rsci_vd),
      .d(chn_o_rsci_d),
      .lz(chn_o_rsc_lz),
      .vz(chn_o_rsc_vz),
      .z(chn_o_rsc_z)
    );
  HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_ctrl HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_ld_core_psct(chn_o_rsci_ld_core_psct),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt),
      .chn_o_rsci_ld_core_sct(chn_o_rsci_ld_core_sct),
      .chn_o_rsci_vd(chn_o_rsci_vd)
    );
  HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_dp HLS_fp32_mul_core_chn_o_rsci_chn_o_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_b_rsci
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_b_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsc_z, chn_b_rsc_vz, chn_b_rsc_lz, chn_b_rsci_oswt,
      core_wen, core_wten, chn_b_rsci_iswt0, chn_b_rsci_bawt, chn_b_rsci_wen_comp,
      chn_b_rsci_ld_core_psct, chn_b_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  input chn_b_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_b_rsci_iswt0;
  output chn_b_rsci_bawt;
  output chn_b_rsci_wen_comp;
  input chn_b_rsci_ld_core_psct;
  output [31:0] chn_b_rsci_d_mxwt;


  // Interconnect Declarations
  wire chn_b_rsci_biwt;
  wire chn_b_rsci_bdwt;
  wire chn_b_rsci_ld_core_sct;
  wire chn_b_rsci_vd;
  wire [31:0] chn_b_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP32_MUL_mgc_in_wire_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) chn_b_rsci (
      .ld(chn_b_rsci_ld_core_sct),
      .vd(chn_b_rsci_vd),
      .d(chn_b_rsci_d),
      .lz(chn_b_rsc_lz),
      .vz(chn_b_rsc_vz),
      .z(chn_b_rsc_z)
    );
  HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_ctrl HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_b_rsci_iswt0(chn_b_rsci_iswt0),
      .chn_b_rsci_ld_core_psct(chn_b_rsci_ld_core_psct),
      .chn_b_rsci_biwt(chn_b_rsci_biwt),
      .chn_b_rsci_bdwt(chn_b_rsci_bdwt),
      .chn_b_rsci_ld_core_sct(chn_b_rsci_ld_core_sct),
      .chn_b_rsci_vd(chn_b_rsci_vd)
    );
  HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_dp HLS_fp32_mul_core_chn_b_rsci_chn_b_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .chn_b_rsci_bawt(chn_b_rsci_bawt),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_b_rsci_d_mxwt(chn_b_rsci_d_mxwt),
      .chn_b_rsci_biwt(chn_b_rsci_biwt),
      .chn_b_rsci_bdwt(chn_b_rsci_bdwt),
      .chn_b_rsci_d(chn_b_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core_chn_a_rsci
// ------------------------------------------------------------------


module HLS_fp32_mul_core_chn_a_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_a_rsci_oswt,
      core_wen, chn_a_rsci_iswt0, chn_a_rsci_bawt, chn_a_rsci_wen_comp, chn_a_rsci_ld_core_psct,
      chn_a_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  input chn_a_rsci_ld_core_psct;
  output [31:0] chn_a_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_a_rsci_biwt;
  wire chn_a_rsci_bdwt;
  wire chn_a_rsci_ld_core_sct;
  wire chn_a_rsci_vd;
  wire [31:0] chn_a_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP32_MUL_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd32)) chn_a_rsci (
      .ld(chn_a_rsci_ld_core_sct),
      .vd(chn_a_rsci_vd),
      .d(chn_a_rsci_d),
      .lz(chn_a_rsc_lz),
      .vz(chn_a_rsc_vz),
      .z(chn_a_rsc_z)
    );
  HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_ctrl HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_ld_core_sct(chn_a_rsci_ld_core_sct),
      .chn_a_rsci_vd(chn_a_rsci_vd)
    );
  HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_dp HLS_fp32_mul_core_chn_a_rsci_chn_a_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_d(chn_a_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul_core
// ------------------------------------------------------------------


module HLS_fp32_mul_core (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_b_rsc_z,
      chn_b_rsc_vz, chn_b_rsc_lz, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_a_rsci_oswt,
      chn_b_rsci_oswt, chn_o_rsci_oswt, chn_o_rsci_oswt_unreg, chn_a_rsci_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input [31:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  output [31:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_a_rsci_oswt;
  input chn_b_rsci_oswt;
  input chn_o_rsci_oswt;
  output chn_o_rsci_oswt_unreg;
  output chn_a_rsci_oswt_unreg_pff;


  // Interconnect Declarations
  wire core_wen;
  wire chn_a_rsci_bawt;
  wire chn_a_rsci_wen_comp;
  wire [31:0] chn_a_rsci_d_mxwt;
  wire core_wten;
  wire chn_b_rsci_bawt;
  wire chn_b_rsci_wen_comp;
  wire [31:0] chn_b_rsci_d_mxwt;
  reg chn_o_rsci_iswt0;
  wire chn_o_rsci_bawt;
  wire chn_o_rsci_wen_comp;
  reg chn_o_rsci_d_31;
  reg [7:0] chn_o_rsci_d_30_23;
  reg [22:0] chn_o_rsci_d_22_0;
  wire [1:0] fsm_output;
  wire IsNaN_8U_23U_nor_tmp;
  wire FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp;
  wire [47:0] FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire IsNaN_8U_23U_1_nor_tmp;
  wire mux_tmp;
  wire mux_tmp_1;
  wire or_tmp_24;
  wire mux_tmp_4;
  wire not_tmp_9;
  wire or_tmp_32;
  wire mux_tmp_9;
  wire mux_tmp_10;
  wire or_tmp_36;
  wire mux_tmp_14;
  wire or_tmp_51;
  wire and_dcpl_3;
  wire and_dcpl_6;
  wire and_dcpl_12;
  wire and_dcpl_13;
  wire and_dcpl_16;
  wire and_dcpl_26;
  wire or_tmp_55;
  wire or_tmp_59;
  wire or_tmp_65;
  reg FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_sva;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_3;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_4;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_3;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_4;
  reg FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg [47:0] FpMul_8U_23U_p_mant_p1_sva_2;
  reg [7:0] FpMul_8U_23U_p_expo_sva_5;
  wire [8:0] nl_FpMul_8U_23U_p_expo_sva_5;
  reg IsNaN_8U_23U_land_lpi_1_dfm_4;
  reg [7:0] FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_acc_1_sdt_8_1_itm_2;
  reg [7:0] FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_30_23_itm_2;
  reg FpMul_8U_23U_mux_10_itm_3;
  reg FpMul_8U_23U_mux_10_itm_4;
  reg [22:0] FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_22_0_itm_2;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  reg FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_2;
  reg FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_3;
  reg [30:0] FpMul_8U_23U_ua_sva_1_30_0_1;
  reg [30:0] FpMul_8U_23U_ub_sva_1_30_0_1;
  wire main_stage_en_1;
  wire FpMantRNE_48U_24U_else_and_svs;
  wire FpMul_8U_23U_is_inf_lpi_1_dfm_2;
  wire FpMantRNE_48U_24U_else_carry_sva;
  wire [7:0] FpMul_8U_23U_o_expo_lpi_1_dfm;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0;
  reg reg_chn_b_rsci_iswt0_cse;
  reg reg_chn_b_rsci_ld_core_psct_cse;
  wire chn_o_and_cse;
  reg reg_chn_o_rsci_ld_core_psct_cse;
  wire or_10_cse;
  wire nand_8_cse;
  wire nand_cse;
  wire or_45_cse;
  wire FpMul_8U_23U_or_2_cse;
  wire nor_4_cse;
  wire and_cse;
  wire or_65_cse;
  wire or_29_cse;
  wire mux_24_cse;
  wire and_41_rgt;
  wire and_45_rgt;
  wire and_54_rgt;
  wire and_64_rgt;
  wire and_65_rgt;
  wire mux_20_itm;
  wire chn_o_rsci_d_30_23_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire [7:0] FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0;
  wire FpMul_8U_23U_lor_2_lpi_1_dfm;
  wire IsNaN_8U_23U_aelse_and_cse;
  wire IsNaN_8U_23U_1_aelse_and_cse;
  wire FpMul_8U_23U_ub_FpBitsToFloat_8U_23U_1_or_1_cse;
  wire FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;

  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_1_nl;
  wire[22:0] FpMul_8U_23U_nor_nl;
  wire[22:0] mux_34_nl;
  wire[22:0] FpMantRNE_48U_24U_else_acc_nl;
  wire[23:0] nl_FpMantRNE_48U_24U_else_acc_nl;
  wire[0:0] or_nl;
  wire[7:0] FpMul_8U_23U_FpMul_8U_23U_and_2_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_1_nl;
  wire[0:0] FpBitsToFloat_8U_23U_1_and_nl;
  wire[8:0] FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_FpMul_8U_23U_else_2_acc_1_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_2_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_2_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] nor_32_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] or_25_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] or_33_nl;
  wire[0:0] and_10_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] and_11_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] and_93_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] and_90_nl;
  wire[0:0] FpMul_8U_23U_xor_1_nl;
  wire[0:0] and_95_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] and_91_nl;
  wire[0:0] nand_6_nl;
  wire[8:0] FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_1_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_1_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] asn_FpMul_8U_23U_p_expo_lpi_1_dfm_1_FpMul_8U_23U_else_2_else_and_nl;
  wire[0:0] FpMul_8U_23U_FpMul_8U_23U_nor_1_nl;
  wire[0:0] FpMul_8U_23U_or_1_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl;
  wire[0:0] or_3_nl;
  wire[0:0] nor_nl;
  wire[0:0] or_1_nl;
  wire[0:0] or_7_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] or_22_nl;
  wire[0:0] nor_22_nl;
  wire[0:0] or_39_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_HLS_fp32_mul_core_chn_o_rsci_inst_chn_o_rsci_d;
  assign nl_HLS_fp32_mul_core_chn_o_rsci_inst_chn_o_rsci_d = {chn_o_rsci_d_31 , chn_o_rsci_d_30_23
      , chn_o_rsci_d_22_0};
  HLS_fp32_mul_core_chn_a_rsci HLS_fp32_mul_core_chn_a_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(reg_chn_b_rsci_iswt0_cse),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_ld_core_psct(reg_chn_b_rsci_ld_core_psct_cse),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  HLS_fp32_mul_core_chn_b_rsci HLS_fp32_mul_core_chn_b_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsc_z(chn_b_rsc_z),
      .chn_b_rsc_vz(chn_b_rsc_vz),
      .chn_b_rsc_lz(chn_b_rsc_lz),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_b_rsci_iswt0(reg_chn_b_rsci_iswt0_cse),
      .chn_b_rsci_bawt(chn_b_rsci_bawt),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_b_rsci_ld_core_psct(reg_chn_b_rsci_ld_core_psct_cse),
      .chn_b_rsci_d_mxwt(chn_b_rsci_d_mxwt)
    );
  HLS_fp32_mul_core_chn_o_rsci HLS_fp32_mul_core_chn_o_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_ld_core_psct(reg_chn_o_rsci_ld_core_psct_cse),
      .chn_o_rsci_d(nl_HLS_fp32_mul_core_chn_o_rsci_inst_chn_o_rsci_d[31:0])
    );
  HLS_fp32_mul_core_staller HLS_fp32_mul_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp)
    );
  HLS_fp32_mul_core_core_fsm HLS_fp32_mul_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign iMantWidth_oMantWidth_prb = MUX_s_1_2_2((MUX1HOT_s_1_1_2(1'b1, fsm_output[0])),
      (MUX1HOT_s_1_1_2(1'b1, main_stage_en_1 & (fsm_output[1]))), fsm_output[1]);
  // assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 386
  // PSL HLS_fp32_mul_core_nvdla_float_h_ln386_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign chn_o_and_cse = core_wen & (~(and_dcpl_6 | (~ main_stage_v_2)));
  assign FpMul_8U_23U_or_2_cse = IsNaN_8U_23U_1_land_lpi_1_dfm_4 | IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign IsNaN_8U_23U_aelse_and_cse = core_wen & (~ and_dcpl_6) & mux_tmp_1;
  assign or_10_cse = (~ reg_chn_o_rsci_ld_core_psct_cse) | chn_o_rsci_bawt;
  assign and_41_rgt = or_10_cse & or_29_cse;
  assign or_29_cse = (~ FpMul_8U_23U_else_2_if_acc_itm_8_1) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign nor_4_cse = ~(IsNaN_8U_23U_land_lpi_1_dfm_st_3 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_3));
  assign FpMul_8U_23U_ub_FpBitsToFloat_8U_23U_1_or_1_cse = (or_10_cse & (~ IsNaN_8U_23U_land_lpi_1_dfm_st_3))
      | and_dcpl_26;
  assign IsNaN_8U_23U_1_aelse_and_cse = core_wen & (~ and_dcpl_6) & mux_tmp_4;
  assign and_45_rgt = or_10_cse & FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign or_65_cse = (~ main_stage_v_1) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign nand_8_cse = ~((chn_b_rsci_d_mxwt[30:23]==8'b11111111));
  assign nand_cse = ~((chn_a_rsci_d_mxwt[30:23]==8'b11111111));
  assign and_54_rgt = or_10_cse & (chn_a_rsci_d_mxwt[30:23]==8'b11111111) & (~ IsNaN_8U_23U_nor_tmp);
  assign and_64_rgt = ((chn_a_rsci_d_mxwt[30:23]!=8'b11111111) | IsNaN_8U_23U_nor_tmp)
      & (chn_b_rsci_d_mxwt[30:23]==8'b11111111) & (~ IsNaN_8U_23U_1_nor_tmp) & or_10_cse;
  assign and_90_nl = nand_cse & or_tmp_55;
  assign mux_33_nl = MUX_s_1_2_2((and_90_nl), or_tmp_55, IsNaN_8U_23U_nor_tmp);
  assign and_65_rgt = (mux_33_nl) & or_10_cse;
  assign or_45_cse = FpMul_8U_23U_oelse_1_acc_itm_9_1 | FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp;
  assign and_95_nl = nand_cse & and_cse;
  assign mux_24_cse = MUX_s_1_2_2((and_95_nl), and_cse, IsNaN_8U_23U_nor_tmp);
  assign IsNaN_8U_23U_nor_tmp = ~((chn_a_rsci_d_mxwt[22:0]!=23'b00000000000000000000000));
  assign FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({1'b1 , (FpMul_8U_23U_ua_sva_1_30_0_1[22:0])})
      * ({1'b1 , (FpMul_8U_23U_ub_sva_1_30_0_1[22:0])}));
  assign nl_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_acc_1_sdt_8_1_itm_2)
      + 9'b101000001;
  assign FpMul_8U_23U_else_2_if_acc_nl = nl_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((FpMul_8U_23U_else_2_if_acc_nl));
  assign IsNaN_8U_23U_1_nor_tmp = ~((chn_b_rsci_d_mxwt[22:0]!=23'b00000000000000000000000));
  assign nl_FpMul_8U_23U_oelse_1_acc_1_nl = conv_u2s_8_9(chn_b_rsci_d_mxwt[30:23])
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_1_nl = nl_FpMul_8U_23U_oelse_1_acc_1_nl[8:0];
  assign nl_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_1_nl)
      + conv_u2s_8_10(chn_a_rsci_d_mxwt[30:23]);
  assign FpMul_8U_23U_oelse_1_acc_nl = nl_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((FpMul_8U_23U_oelse_1_acc_nl));
  assign FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp = (~((chn_b_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000)))
      | (~((chn_a_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000)));
  assign nl_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_sva_5[7:1])})
      + 8'b1;
  assign FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = readslicef_8_1_7((FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign nl_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_sva_5 + 8'b1;
  assign FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign asn_FpMul_8U_23U_p_expo_lpi_1_dfm_1_FpMul_8U_23U_else_2_else_and_nl = FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      & (FpMul_8U_23U_p_mant_p1_sva_2[47]);
  assign FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0 = MUX_v_8_2_2(FpMul_8U_23U_p_expo_sva_5,
      (FpMul_8U_23U_else_2_else_if_if_acc_nl), asn_FpMul_8U_23U_p_expo_lpi_1_dfm_1_FpMul_8U_23U_else_2_else_and_nl);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1[7:0];
  assign FpMantRNE_48U_24U_else_and_svs = FpMantRNE_48U_24U_else_carry_sva & (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_sva = (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_sva_2[0]) & (FpMul_8U_23U_p_mant_p1_sva_2[47]))
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_sva_2[45:0]),
      (FpMul_8U_23U_p_mant_p1_sva_2[46:1]), FpMul_8U_23U_p_mant_p1_sva_2[47]);
  assign FpMul_8U_23U_FpMul_8U_23U_nor_1_nl = ~(FpMantRNE_48U_24U_else_and_svs |
      FpMul_8U_23U_is_inf_lpi_1_dfm_2);
  assign FpMul_8U_23U_or_1_nl = ((~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp)
      & FpMantRNE_48U_24U_else_and_svs) | FpMul_8U_23U_is_inf_lpi_1_dfm_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp
      & FpMantRNE_48U_24U_else_and_svs & (~ FpMul_8U_23U_is_inf_lpi_1_dfm_2);
  assign FpMul_8U_23U_o_expo_lpi_1_dfm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1, {(FpMul_8U_23U_FpMul_8U_23U_nor_1_nl)
      , (FpMul_8U_23U_or_1_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl)});
  assign FpMul_8U_23U_lor_2_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_lpi_1_dfm!=8'b00000000)))
      | FpMul_8U_23U_lor_1_lpi_1_dfm_4;
  assign FpMul_8U_23U_is_inf_lpi_1_dfm_2 = ~(((FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | (~ (FpMul_8U_23U_p_mant_p1_sva_2[47]))) & FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_4);
  assign main_stage_en_1 = chn_a_rsci_bawt & chn_b_rsci_bawt & or_10_cse;
  assign or_3_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ main_stage_v_1) | chn_o_rsci_bawt
      | (~ reg_chn_o_rsci_ld_core_psct_cse);
  assign nor_nl = ~((~(FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ main_stage_v_1))) |
      chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign or_1_nl = (~ chn_a_rsci_bawt) | (~ chn_b_rsci_bawt) | FpMul_8U_23U_oelse_1_acc_itm_9_1
      | FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp;
  assign mux_tmp = MUX_s_1_2_2((nor_nl), (or_3_nl), or_1_nl);
  assign and_cse = chn_a_rsci_bawt & chn_b_rsci_bawt;
  assign or_7_nl = main_stage_v_1 | chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse);
  assign nor_28_nl = ~((~ main_stage_v_1) | chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign mux_tmp_1 = MUX_s_1_2_2((nor_28_nl), (or_7_nl), and_cse);
  assign or_tmp_24 = (~ main_stage_v_2) | chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse);
  assign or_22_nl = main_stage_v_2 | chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse);
  assign mux_tmp_4 = MUX_s_1_2_2((~ or_tmp_24), (or_22_nl), main_stage_v_1);
  assign not_tmp_9 = ~(main_stage_v_1 & or_10_cse);
  assign or_tmp_32 = (~(chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse))) |
      IsNaN_8U_23U_land_lpi_1_dfm_st_3;
  assign nor_22_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ IsNaN_8U_23U_land_lpi_1_dfm_st_3));
  assign mux_tmp_9 = MUX_s_1_2_2((nor_22_nl), IsNaN_8U_23U_land_lpi_1_dfm_st_3, chn_o_rsci_bawt);
  assign mux_tmp_10 = MUX_s_1_2_2(mux_tmp_9, or_10_cse, nor_4_cse);
  assign or_tmp_36 = IsNaN_8U_23U_1_land_lpi_1_dfm_3 | or_tmp_32;
  assign mux_tmp_14 = MUX_s_1_2_2(mux_tmp_9, or_10_cse, IsNaN_8U_23U_1_land_lpi_1_dfm_3);
  assign or_39_nl = (~ main_stage_v_1) | IsNaN_8U_23U_1_land_lpi_1_dfm_3 | or_tmp_32;
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_36, mux_tmp_14, main_stage_v_2);
  assign mux_19_nl = MUX_s_1_2_2(or_tmp_24, (mux_18_nl), main_stage_v_1);
  assign mux_20_itm = MUX_s_1_2_2((mux_19_nl), (or_39_nl), FpMul_8U_23U_or_2_cse);
  assign or_tmp_51 = FpMul_8U_23U_oelse_1_acc_itm_9_1 | FpMul_8U_23U_if_2_FpMul_8U_23U_if_2_or_tmp
      | (~ and_cse);
  assign and_dcpl_3 = chn_o_rsci_bawt & reg_chn_o_rsci_ld_core_psct_cse;
  assign and_dcpl_6 = (~ chn_o_rsci_bawt) & reg_chn_o_rsci_ld_core_psct_cse;
  assign and_dcpl_12 = or_10_cse & main_stage_v_2;
  assign and_dcpl_13 = and_dcpl_3 & (~ main_stage_v_2);
  assign and_dcpl_16 = or_10_cse & main_stage_v_1;
  assign and_dcpl_26 = or_10_cse & IsNaN_8U_23U_land_lpi_1_dfm_st_3;
  assign or_tmp_55 = IsNaN_8U_23U_1_nor_tmp | nand_8_cse;
  assign or_tmp_59 = main_stage_en_1 | (fsm_output[0]);
  assign or_tmp_65 = or_10_cse & chn_b_rsci_bawt & chn_a_rsci_bawt & (fsm_output[1]);
  assign chn_o_rsci_d_30_23_mx0c1 = or_10_cse & main_stage_v_2 & (~ IsNaN_8U_23U_land_lpi_1_dfm_4);
  assign main_stage_v_1_mx0c1 = and_dcpl_16 & (~(chn_b_rsci_bawt & chn_a_rsci_bawt));
  assign main_stage_v_2_mx0c1 = or_10_cse & main_stage_v_2 & (~ main_stage_v_1);
  assign chn_a_rsci_oswt_unreg_pff = or_tmp_65;
  assign chn_o_rsci_oswt_unreg = and_dcpl_3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_b_rsci_iswt0_cse <= 1'b0;
      chn_o_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_chn_b_rsci_iswt0_cse <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_o_rsci_iswt0 <= and_dcpl_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_b_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & or_tmp_59 ) begin
      reg_chn_b_rsci_ld_core_psct_cse <= or_tmp_59;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_22_0 <= 23'b0;
      chn_o_rsci_d_31 <= 1'b0;
    end
    else if ( chn_o_and_cse ) begin
      chn_o_rsci_d_22_0 <= MUX_v_23_2_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_1_nl),
          FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_22_0_itm_2, FpMul_8U_23U_or_2_cse);
      chn_o_rsci_d_31 <= FpMul_8U_23U_mux_10_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_30_23 <= 8'b0;
    end
    else if ( core_wen & ((or_10_cse & main_stage_v_2 & IsNaN_8U_23U_land_lpi_1_dfm_4)
        | chn_o_rsci_d_30_23_mx0c1) ) begin
      chn_o_rsci_d_30_23 <= MUX_v_8_2_2(FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_30_23_itm_2,
          (FpMul_8U_23U_FpMul_8U_23U_and_2_nl), FpBitsToFloat_8U_23U_1_and_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_12 | and_dcpl_13) ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= ~ and_dcpl_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_65 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_acc_1_sdt_8_1_itm_2 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (~ mux_tmp) ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_acc_1_sdt_8_1_itm_2 <= readslicef_9_8_1((FpMul_8U_23U_else_2_acc_1_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_3 <= 1'b0;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_8U_23U_1_land_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_3 <= ~(IsNaN_8U_23U_nor_tmp | nand_cse);
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= or_45_cse;
      IsNaN_8U_23U_1_land_lpi_1_dfm_3 <= ~(IsNaN_8U_23U_1_nor_tmp | nand_8_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_16 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_sva_5 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (mux_3_nl) ) begin
      FpMul_8U_23U_p_expo_sva_5 <= nl_FpMul_8U_23U_p_expo_sva_5[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_sva_2 <= 48'b0;
    end
    else if ( core_wen & ((or_10_cse & (~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_3) & FpMul_8U_23U_else_2_if_acc_itm_8_1)
        | and_41_rgt) & mux_tmp_4 ) begin
      FpMul_8U_23U_p_mant_p1_sva_2 <= MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_mul_tmp,
          FpMul_8U_23U_p_mant_p1_sva, and_41_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (mux_6_nl) ) begin
      FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (mux_8_nl) ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_2 <= FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_30_23_itm_2 <= 8'b0;
    end
    else if ( core_wen & FpMul_8U_23U_ub_FpBitsToFloat_8U_23U_1_or_1_cse & (mux_13_nl)
        ) begin
      FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_30_23_itm_2 <= MUX_v_8_2_2((FpMul_8U_23U_ub_sva_1_30_0_1[30:23]),
          (FpMul_8U_23U_ua_sva_1_30_0_1[30:23]), and_dcpl_26);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_4 <= 1'b0;
      FpMul_8U_23U_mux_10_itm_4 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_cse ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_4 <= IsNaN_8U_23U_1_land_lpi_1_dfm_3;
      FpMul_8U_23U_mux_10_itm_4 <= FpMul_8U_23U_mux_10_itm_3;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= IsNaN_8U_23U_land_lpi_1_dfm_st_3;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_22_0_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpMul_8U_23U_ub_FpBitsToFloat_8U_23U_1_or_1_cse & (mux_17_nl)
        ) begin
      FpBitsToFloat_8U_23U_1_slc_FpBitsToFloat_8U_23U_ubits_1_22_0_itm_2 <= MUX_v_23_2_2((FpMul_8U_23U_ub_sva_1_30_0_1[22:0]),
          (FpMul_8U_23U_ua_sva_1_30_0_1[22:0]), and_dcpl_26);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (~ mux_20_itm) ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_4 <= FpMul_8U_23U_lor_1_lpi_1_dfm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_10_cse & (~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_3)) | and_45_rgt)
        & (~ mux_20_itm) ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_if_acc_itm_8_1,
          FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs, and_45_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_sva <= 48'b0;
    end
    else if ( core_wen & (~(and_dcpl_6 | (~ main_stage_v_1) | or_29_cse)) ) begin
      FpMul_8U_23U_p_mant_p1_sva <= FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~ (fsm_output[0])) & (~ or_65_cse) & mux_tmp ) begin
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (mux_23_nl) ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_3 <= or_45_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_10_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_54_rgt | and_64_rgt | and_65_rgt) & mux_tmp_1 ) begin
      FpMul_8U_23U_mux_10_itm_3 <= MUX1HOT_s_1_3_2((chn_a_rsci_d_mxwt[31]), (chn_b_rsci_d_mxwt[31]),
          (FpMul_8U_23U_xor_1_nl), {and_54_rgt , and_64_rgt , and_65_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_ub_sva_1_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (mux_28_nl) ) begin
      FpMul_8U_23U_ub_sva_1_30_0_1 <= chn_b_rsci_d_mxwt[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_ua_sva_1_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_6) & (~ (mux_31_nl)) ) begin
      FpMul_8U_23U_ua_sva_1_30_0_1 <= chn_a_rsci_d_mxwt[30:0];
    end
  end
  assign nl_FpMantRNE_48U_24U_else_acc_nl = (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23])
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_sva);
  assign FpMantRNE_48U_24U_else_acc_nl = nl_FpMantRNE_48U_24U_else_acc_nl[22:0];
  assign or_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp | (~ FpMantRNE_48U_24U_else_and_svs);
  assign mux_34_nl = MUX_v_23_2_2((signext_23_1(~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp)),
      (FpMantRNE_48U_24U_else_acc_nl), or_nl);
  assign FpMul_8U_23U_nor_nl = ~(MUX_v_23_2_2((mux_34_nl), 23'b11111111111111111111111,
      FpMul_8U_23U_is_inf_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_1_nl = ~(MUX_v_23_2_2((FpMul_8U_23U_nor_nl),
      23'b11111111111111111111111, FpMul_8U_23U_lor_2_lpi_1_dfm));
  assign FpMul_8U_23U_oelse_2_not_1_nl = ~ FpMul_8U_23U_lor_2_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_2_nl = MUX_v_8_2_2(8'b00000000, FpMul_8U_23U_o_expo_lpi_1_dfm,
      (FpMul_8U_23U_oelse_2_not_1_nl));
  assign FpBitsToFloat_8U_23U_1_and_nl = (~ IsNaN_8U_23U_1_land_lpi_1_dfm_4) & chn_o_rsci_d_30_23_mx0c1;
  assign nl_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(chn_a_rsci_d_mxwt[30:23])
      + conv_u2u_8_9(chn_b_rsci_d_mxwt[30:23]);
  assign FpMul_8U_23U_else_2_acc_1_nl = nl_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_FpMul_8U_23U_else_2_else_acc_2_nl = (FpMul_8U_23U_ub_sva_1_30_0_1[30:23])
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_2_nl = nl_FpMul_8U_23U_else_2_else_acc_2_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_sva_5  = (FpMul_8U_23U_else_2_else_acc_2_nl) + (FpMul_8U_23U_ua_sva_1_30_0_1[30:23]);
  assign nor_24_nl = ~((~ main_stage_v_1) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~(FpMul_8U_23U_else_2_if_acc_itm_8_1
      & ((FpMul_8U_23U_p_mant_p1_mul_tmp[47]) | (~(IsNaN_8U_23U_land_lpi_1_dfm_st_3
      | IsNaN_8U_23U_1_land_lpi_1_dfm_3))))));
  assign nor_26_nl = ~((~ main_stage_v_2) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | (~
      FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_2));
  assign nor_27_nl = ~(FpMul_8U_23U_or_2_cse | (FpMul_8U_23U_p_mant_p1_sva_2[47])
      | (~ main_stage_v_2) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | (~ FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_2));
  assign mux_2_nl = MUX_s_1_2_2((nor_27_nl), (nor_26_nl), FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2);
  assign mux_3_nl = MUX_s_1_2_2((mux_2_nl), (nor_24_nl), or_10_cse);
  assign nor_32_nl = ~((~ FpMul_8U_23U_else_2_if_acc_itm_8_1) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | not_tmp_9);
  assign mux_5_nl = MUX_s_1_2_2(mux_tmp_4, (~ or_tmp_24), or_29_cse);
  assign or_25_nl = (~ FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_2)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  assign mux_6_nl = MUX_s_1_2_2((mux_5_nl), (nor_32_nl), or_25_nl);
  assign nor_23_nl = ~(FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | not_tmp_9);
  assign mux_7_nl = MUX_s_1_2_2(mux_tmp_4, (~ or_tmp_24), FpMul_8U_23U_lor_1_lpi_1_dfm_st_3);
  assign mux_8_nl = MUX_s_1_2_2((mux_7_nl), (nor_23_nl), FpMul_8U_23U_lor_1_lpi_1_dfm_st_4);
  assign or_33_nl = nor_4_cse | or_tmp_32;
  assign mux_11_nl = MUX_s_1_2_2(mux_tmp_10, (or_33_nl), main_stage_v_2);
  assign mux_12_nl = MUX_s_1_2_2((~ or_tmp_24), (mux_11_nl), main_stage_v_1);
  assign and_10_nl = main_stage_v_1 & mux_tmp_10;
  assign mux_13_nl = MUX_s_1_2_2((and_10_nl), (mux_12_nl), FpMul_8U_23U_or_2_cse);
  assign mux_15_nl = MUX_s_1_2_2(mux_tmp_14, or_tmp_36, main_stage_v_2);
  assign mux_16_nl = MUX_s_1_2_2((~ or_tmp_24), (mux_15_nl), main_stage_v_1);
  assign and_11_nl = main_stage_v_1 & mux_tmp_14;
  assign mux_17_nl = MUX_s_1_2_2((and_11_nl), (mux_16_nl), FpMul_8U_23U_or_2_cse);
  assign and_93_nl = nand_8_cse & mux_24_cse;
  assign mux_22_nl = MUX_s_1_2_2((and_93_nl), mux_24_cse, IsNaN_8U_23U_1_nor_tmp);
  assign nor_21_nl = ~((~ main_stage_v_1) | IsNaN_8U_23U_land_lpi_1_dfm_st_3 | IsNaN_8U_23U_1_land_lpi_1_dfm_3);
  assign mux_23_nl = MUX_s_1_2_2((nor_21_nl), (mux_22_nl), or_10_cse);
  assign FpMul_8U_23U_xor_1_nl = (chn_a_rsci_d_mxwt[31]) ^ (chn_b_rsci_d_mxwt[31]);
  assign nor_31_nl = ~(IsNaN_8U_23U_1_nor_tmp | (~((chn_b_rsci_d_mxwt[30:23]==8'b11111111)
      & mux_24_cse)));
  assign mux_25_nl = MUX_s_1_2_2(and_cse, (nor_31_nl), or_45_cse);
  assign mux_26_nl = MUX_s_1_2_2(or_65_cse, (~ main_stage_v_1), IsNaN_8U_23U_1_land_lpi_1_dfm_3);
  assign mux_27_nl = MUX_s_1_2_2((mux_26_nl), or_65_cse, IsNaN_8U_23U_land_lpi_1_dfm_st_3);
  assign mux_28_nl = MUX_s_1_2_2((~ (mux_27_nl)), (mux_25_nl), or_10_cse);
  assign and_91_nl = (chn_a_rsci_d_mxwt[30:23]==8'b11111111);
  assign mux_29_nl = MUX_s_1_2_2(or_tmp_51, (~ and_cse), and_91_nl);
  assign mux_30_nl = MUX_s_1_2_2((mux_29_nl), or_tmp_51, IsNaN_8U_23U_nor_tmp);
  assign nand_6_nl = ~(((~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_3) | IsNaN_8U_23U_land_lpi_1_dfm_st_3)
      & main_stage_v_1);
  assign mux_31_nl = MUX_s_1_2_2((nand_6_nl), (mux_30_nl), or_10_cse);

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [45:0] MUX_v_46_2_2;
    input [45:0] input_0;
    input [45:0] input_1;
    input [0:0] sel;
    reg [45:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_46_2_2 = result;
  end
  endfunction


  function [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function [22:0] signext_23_1;
    input [0:0] vector;
  begin
    signext_23_1= {{22{vector[0]}}, vector};
  end
  endfunction


  function  [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function  [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function  [9:0] conv_u2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [22:0] conv_u2u_1_23 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction


  function  [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function  [47:0] conv_u2u_48_48 ;
    input [47:0]  vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_mul
// ------------------------------------------------------------------


module HLS_fp32_mul (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_b_rsc_z,
      chn_b_rsc_vz, chn_b_rsc_lz, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input [31:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  output [31:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;


  // Interconnect Declarations
  wire chn_a_rsci_oswt;
  wire chn_b_rsci_oswt;
  wire chn_o_rsci_oswt;
  wire chn_o_rsci_oswt_unreg;
  wire chn_a_rsci_oswt_unreg_iff;


  // Interconnect Declarations for Component Instantiations 
  FP32_MUL_chn_a_rsci_unreg chn_a_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg_iff),
      .outsig(chn_a_rsci_oswt)
    );
  FP32_MUL_chn_b_rsci_unreg chn_b_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg_iff),
      .outsig(chn_b_rsci_oswt)
    );
  FP32_MUL_chn_o_rsci_unreg chn_o_rsci_unreg_inst (
      .in_0(chn_o_rsci_oswt_unreg),
      .outsig(chn_o_rsci_oswt)
    );
  HLS_fp32_mul_core HLS_fp32_mul_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_b_rsc_z(chn_b_rsc_z),
      .chn_b_rsc_vz(chn_b_rsc_vz),
      .chn_b_rsc_lz(chn_b_rsc_lz),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_oswt_unreg(chn_o_rsci_oswt_unreg),
      .chn_a_rsci_oswt_unreg_pff(chn_a_rsci_oswt_unreg_iff)
    );
endmodule



