// Common coverage definition

`define PDP_COV_BIN_NUM_DEFAULT         8
`define CDP_COV_BIN_NUM_DEFAULT         8
`define MAX_VALUE_27BITS                27'h7FF_FFFF
`define MAX_VALUE_8BITS                 8'hFF
`define MAX_VALUE_3BITS                 3'h7

