// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// nvdla_top sv side SC-SV Adapter 
// This is autogenerated code 

`ifndef _nvdla_top_sv_tlm_callbacks
`define _nvdla_top_sv_tlm_callbacks

class nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks);

    /// Creates a new nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks
    function new(string name = "nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
        dbb_bus_ext dbb_bus_tr;
        $cast(dbb_bus_tr, obj.get_extension(dbb_bus_ext::ID));
        obj.set_transaction_id(dbb_bus_tr.get_id);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks
                  
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
class nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks);

    /// Creates a new nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks
    function new(string name = "nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
        dbb_bus_ext dbb_bus_tr;
        $cast(dbb_bus_tr, obj.get_extension(dbb_bus_ext::ID));
        obj.set_transaction_id(dbb_bus_tr.get_id);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks
`endif
                  
class nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks);

    /// Creates a new nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks
    function new(string name = "nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks
                  
class nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks);

    /// Creates a new nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks
    function new(string name = "nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks
                  
class nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks);

    /// Creates a new nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks
    function new(string name = "nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks
                  
class nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks);

    /// Creates a new nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks
    function new(string name = "nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks
                  
class nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks);

    /// Creates a new nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks
    function new(string name = "nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks
                  
class nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks);

    /// Creates a new nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks
    function new(string name = "nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks
                  
class nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks);

    /// Creates a new nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks
    function new(string name = "nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks
                  
class nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks);

    /// Creates a new nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks
    function new(string name = "nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks
                  
class nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks #(type T = tlm_generic_payload) extends nvdla_scsv_sv_tlm_callbacks #(T);

    `uvm_object_utils(nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks);

    /// Creates a new nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks
    function new(string name = "nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks");
        super.new(name);
    endfunction: new

    /// Called before a transaction is executed
    virtual task pre_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: pre_btransport_cb

    /// Called after a transaction has been executed
    virtual task post_btransport_cb(nvdla_scsv_sv_tlm_channel#(T) converter, T obj, uvm_tlm_time delay);
	
    endtask: post_btransport_cb

endclass:nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks
 



//Macro containing callback declarations
//If the compile time define NEED_SCSV_SV_CALLBACKS is passed,
//This shall be used as-is in nvdla_top_sv_layer.svh
`define nvdla_top_DEC_MACRO \
                 nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks_inst;  \
               `ifdef NVDLA_SECONDARY_MEMIF_ENABLE \
               nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks_inst;  \
               `endif \
               nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks_inst;  \
               nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks_inst;  \
               nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks_inst;  \
               nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks_inst;  \
               nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks_inst;  \
               nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks_inst;  \
               nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks_inst;  \
               nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks_inst;  \
               nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks_inst;  \
 



//Macro containing callback object construction calls
//If the compile time define NEED_SCSV_SV_CALLBACKS is passed,
//This shall be used as-is in the build_phase of nvdla_top_sv_layer.svh
`define nvdla_top_CONSTRUCT_MACRO \
                 nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks_inst = nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks_inst",this);  \
               `ifdef NVDLA_SECONDARY_MEMIF_ENABLE \
               nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks_inst = nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks_inst",this);  \
               `endif \
               nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks_inst = nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks_inst",this);  \
               nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks_inst = nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks_inst",this);  \
               nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks_inst = nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks_inst",this);  \
               nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks_inst = nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks_inst",this);  \
               nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks_inst = nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks_inst",this);  \
               nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks_inst = nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks_inst",this);  \
               nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks_inst = nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks_inst",this);  \
               nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks_inst = nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks_inst",this);  \
               nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks_inst = nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks_inst",this);  \
 



//Macro containing callback registration calls
//If the compile time define NEED_SCSV_SV_CALLBACKS is passed,
//This shall be used as-is in the connect_phase of nvdla_top_sv_layer.svh
`define nvdla_top_REGISTER_MACRO \
                 uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sc2sv_nvdla_core2dbb_axi4,nvdla_top_sc2sv_nvdla_core2dbb_axi4_tlm_callbacks_inst);  \
               `ifdef NVDLA_SECONDARY_MEMIF_ENABLE \
               uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sc2sv_nvdla_core2cvsram_axi4,nvdla_top_sc2sv_nvdla_core2cvsram_axi4_tlm_callbacks_inst);  \
               `endif \
               uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sv2sc_nvdla_host_master_if,nvdla_top_sv2sc_nvdla_host_master_if_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sc2sv_dma_monitor_mc,nvdla_top_sc2sv_dma_monitor_mc_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sc2sv_dma_monitor_cv,nvdla_top_sc2sv_dma_monitor_cv_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sc2sv_convolution_core_monitor_initiator,nvdla_top_sc2sv_convolution_core_monitor_initiator_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sc2sv_post_processing_monitor_initiator,nvdla_top_sc2sv_post_processing_monitor_initiator_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sv2sc_dma_monitor_mc_credit,nvdla_top_sv2sc_dma_monitor_mc_credit_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sv2sc_dma_monitor_cv_credit,nvdla_top_sv2sc_dma_monitor_cv_credit_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sv2sc_convolution_core_monitor_credit,nvdla_top_sv2sc_convolution_core_monitor_credit_tlm_callbacks_inst);  \
               //uvm_callbacks #(nvdla_scsv_sv_tlm_channel#(tlm_generic_payload), nvdla_scsv_sv_tlm_callbacks#(tlm_generic_payload))::add(nvdla_top_sv2sc_post_processing_monitor_credit,nvdla_top_sv2sc_post_processing_monitor_credit_tlm_callbacks_inst);  \
 


`endif // nvdla_top_sv_tlm_callbacks 
