// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: HLS_fp17_to_fp32.v

module FP17_TO_FP32_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/FP17_TO_FP32_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module FP17_TO_FP32_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-084
//  Generated date: Mon Mar 20 14:09:21 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    FP17_TO_FP32_chn_o_rsci_unreg
// ------------------------------------------------------------------


module FP17_TO_FP32_chn_o_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP17_TO_FP32_chn_a_rsci_unreg
// ------------------------------------------------------------------


module FP17_TO_FP32_chn_a_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for HLS_fp17_to_fp32_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : HLS_fp17_to_fp32_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_staller
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_a_rsci_wen_comp, core_wten, chn_o_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_a_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_o_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_a_rsci_wen_comp & chn_o_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_biwt, chn_o_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_biwt;
  input chn_o_rsci_bdwt;


  // Interconnect Declarations
  reg chn_o_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_bawt = chn_o_rsci_biwt | chn_o_rsci_bcwt;
  assign chn_o_rsci_wen_comp = (~ chn_o_rsci_oswt) | chn_o_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_o_rsci_bcwt <= ~((~(chn_o_rsci_bcwt | chn_o_rsci_biwt)) | chn_o_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, core_wen, core_wten, chn_o_rsci_iswt0,
      chn_o_rsci_ld_core_psct, chn_o_rsci_biwt, chn_o_rsci_bdwt, chn_o_rsci_ld_core_sct,
      chn_o_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  input chn_o_rsci_ld_core_psct;
  output chn_o_rsci_biwt;
  output chn_o_rsci_bdwt;
  output chn_o_rsci_ld_core_sct;
  input chn_o_rsci_vd;


  // Interconnect Declarations
  wire chn_o_rsci_ogwt;
  wire chn_o_rsci_pdswt0;
  reg chn_o_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_pdswt0 = (~ core_wten) & chn_o_rsci_iswt0;
  assign chn_o_rsci_biwt = chn_o_rsci_ogwt & chn_o_rsci_vd;
  assign chn_o_rsci_ogwt = chn_o_rsci_pdswt0 | chn_o_rsci_icwt;
  assign chn_o_rsci_bdwt = chn_o_rsci_oswt & core_wen;
  assign chn_o_rsci_ld_core_sct = chn_o_rsci_ld_core_psct & chn_o_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_icwt <= 1'b0;
    end
    else begin
      chn_o_rsci_icwt <= ~((~(chn_o_rsci_icwt | chn_o_rsci_pdswt0)) | chn_o_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, chn_a_rsci_bawt, chn_a_rsci_wen_comp,
      chn_a_rsci_d_mxwt, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  output [16:0] chn_a_rsci_d_mxwt;
  input chn_a_rsci_biwt;
  input chn_a_rsci_bdwt;
  input [16:0] chn_a_rsci_d;


  // Interconnect Declarations
  reg chn_a_rsci_bcwt;
  reg [16:0] chn_a_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_bawt = chn_a_rsci_biwt | chn_a_rsci_bcwt;
  assign chn_a_rsci_wen_comp = (~ chn_a_rsci_oswt) | chn_a_rsci_bawt;
  assign chn_a_rsci_d_mxwt = MUX_v_17_2_2(chn_a_rsci_d, chn_a_rsci_d_bfwt, chn_a_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_bcwt <= 1'b0;
      chn_a_rsci_d_bfwt <= 17'b0;
    end
    else begin
      chn_a_rsci_bcwt <= ~((~(chn_a_rsci_bcwt | chn_a_rsci_biwt)) | chn_a_rsci_bdwt);
      chn_a_rsci_d_bfwt <= chn_a_rsci_d_mxwt;
    end
  end

  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct,
      core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  input chn_a_rsci_ld_core_psct;
  input core_wten;
  output chn_a_rsci_biwt;
  output chn_a_rsci_bdwt;
  output chn_a_rsci_ld_core_sct;
  input chn_a_rsci_vd;


  // Interconnect Declarations
  wire chn_a_rsci_ogwt;
  wire chn_a_rsci_pdswt0;
  reg chn_a_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_pdswt0 = (~ core_wten) & chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & chn_a_rsci_vd;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | chn_a_rsci_icwt;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & chn_a_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_icwt <= 1'b0;
    end
    else begin
      chn_a_rsci_icwt <= ~((~(chn_a_rsci_icwt | chn_a_rsci_pdswt0)) | chn_a_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_chn_o_rsci
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_chn_o_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_o_rsci_oswt,
      core_wen, core_wten, chn_o_rsci_iswt0, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_ld_core_psct, chn_o_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [31:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_ld_core_psct;
  input [31:0] chn_o_rsci_d;


  // Interconnect Declarations
  wire chn_o_rsci_biwt;
  wire chn_o_rsci_bdwt;
  wire chn_o_rsci_ld_core_sct;
  wire chn_o_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  FP17_TO_FP32_mgc_out_stdreg_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) chn_o_rsci (
      .ld(chn_o_rsci_ld_core_sct),
      .vd(chn_o_rsci_vd),
      .d(chn_o_rsci_d),
      .lz(chn_o_rsc_lz),
      .vz(chn_o_rsc_vz),
      .z(chn_o_rsc_z)
    );
  HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_ctrl HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_ld_core_psct(chn_o_rsci_ld_core_psct),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt),
      .chn_o_rsci_ld_core_sct(chn_o_rsci_ld_core_sct),
      .chn_o_rsci_vd(chn_o_rsci_vd)
    );
  HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_dp HLS_fp17_to_fp32_core_chn_o_rsci_chn_o_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core_chn_a_rsci
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core_chn_a_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_a_rsci_oswt,
      core_wen, chn_a_rsci_iswt0, chn_a_rsci_bawt, chn_a_rsci_wen_comp, chn_a_rsci_ld_core_psct,
      chn_a_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  input chn_a_rsci_ld_core_psct;
  output [16:0] chn_a_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_a_rsci_biwt;
  wire chn_a_rsci_bdwt;
  wire chn_a_rsci_ld_core_sct;
  wire chn_a_rsci_vd;
  wire [16:0] chn_a_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP17_TO_FP32_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd17)) chn_a_rsci (
      .ld(chn_a_rsci_ld_core_sct),
      .vd(chn_a_rsci_vd),
      .d(chn_a_rsci_d),
      .lz(chn_a_rsc_lz),
      .vz(chn_a_rsc_vz),
      .z(chn_a_rsc_z)
    );
  HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_ctrl HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_ld_core_sct(chn_a_rsci_ld_core_sct),
      .chn_a_rsci_vd(chn_a_rsci_vd)
    );
  HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_dp HLS_fp17_to_fp32_core_chn_a_rsci_chn_a_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_d(chn_a_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32_core
// ------------------------------------------------------------------


module HLS_fp17_to_fp32_core (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_o_rsc_z,
      chn_o_rsc_vz, chn_o_rsc_lz, chn_a_rsci_oswt, chn_a_rsci_oswt_unreg, chn_o_rsci_oswt,
      chn_o_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  output [31:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_a_rsci_oswt;
  output chn_a_rsci_oswt_unreg;
  input chn_o_rsci_oswt;
  output chn_o_rsci_oswt_unreg;


  // Interconnect Declarations
  wire core_wen;
  reg chn_a_rsci_iswt0;
  wire chn_a_rsci_bawt;
  wire chn_a_rsci_wen_comp;
  reg chn_a_rsci_ld_core_psct;
  wire [16:0] chn_a_rsci_d_mxwt;
  wire core_wten;
  wire chn_o_rsci_bawt;
  wire chn_o_rsci_wen_comp;
  reg chn_o_rsci_d_31;
  reg [2:0] chn_o_rsci_d_30_28;
  reg [4:0] chn_o_rsci_d_27_23;
  reg [9:0] chn_o_rsci_d_22_13;
  reg [9:0] chn_o_rsci_d_9_0;
  reg chn_o_rsci_d_10;
  wire [1:0] fsm_output;
  wire IsNaN_6U_23U_nor_tmp;
  wire and_dcpl_2;
  wire or_dcpl_3;
  wire and_dcpl_7;
  wire and_dcpl_11;
  wire or_dcpl_9;
  wire and_dcpl_25;
  wire or_tmp_18;
  wire and_46_cse;
  wire and_48_cse;
  wire and_4_mdf;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nand_cse;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm;
  wire chn_o_and_4_cse;
  reg reg_chn_o_rsci_iswt0_cse;
  reg reg_chn_o_rsci_ld_core_psct_cse;
  wire or_cse;
  wire chn_o_rsci_d_9_0_mx0c1;
  wire IsInf_6U_23U_land_lpi_1_dfm_mx1w0;
  wire HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_sig_mx0;
  wire chn_a_rsci_ld_core_psct_mx0c0;
  wire IsNaN_6U_23U_land_lpi_1_dfm;

  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_1;
  wire[0:0] nand_11_nl;
  wire[0:0] nand_10_nl;
  wire[4:0] FpExpoWidthInc_6U_8U_23U_0U_1U_mux_5_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[3:0] nl_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[0:0] IsZero_6U_23U_aelse_IsZero_6U_23U_or_nl;
  wire[0:0] and_6_nl;
  wire[0:0] IsNaN_6U_23U_aelse_not_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_HLS_fp17_to_fp32_core_chn_o_rsci_inst_chn_o_rsci_d;
  assign nl_HLS_fp17_to_fp32_core_chn_o_rsci_inst_chn_o_rsci_d = {chn_o_rsci_d_31
      , chn_o_rsci_d_30_28 , chn_o_rsci_d_27_23 , chn_o_rsci_d_22_13 , ({{2{chn_o_rsci_d_10}},
      chn_o_rsci_d_10}) , chn_o_rsci_d_9_0};
  HLS_fp17_to_fp32_core_chn_a_rsci HLS_fp17_to_fp32_core_chn_a_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  HLS_fp17_to_fp32_core_chn_o_rsci HLS_fp17_to_fp32_core_chn_o_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(reg_chn_o_rsci_iswt0_cse),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_ld_core_psct(reg_chn_o_rsci_ld_core_psct_cse),
      .chn_o_rsci_d(nl_HLS_fp17_to_fp32_core_chn_o_rsci_inst_chn_o_rsci_d[31:0])
    );
  HLS_fp17_to_fp32_core_staller HLS_fp17_to_fp32_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp)
    );
  HLS_fp17_to_fp32_core_core_fsm HLS_fp17_to_fp32_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign iExpoWidth_oExpoWidth_prb = HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_sig_mx0;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 596
  // PSL HLS_fp17_to_fp32_core_nvdla_float_h_ln596_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb = HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_sig_mx0;
  // assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 597
  // PSL HLS_fp17_to_fp32_core_nvdla_float_h_ln597_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_1 = HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_sig_mx0;
  // assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 550
  // PSL HLS_fp17_to_fp32_core_nvdla_float_h_ln550_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_1 = HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_sig_mx0;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_1 } @rose(nvdla_core_clk);
  assign chn_o_and_4_cse = core_wen & (~(or_dcpl_3 | (fsm_output[0])));
  assign and_6_nl = and_4_mdf & (fsm_output[1]);
  assign HLS_fp17_to_fp32_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_sig_mx0
      = MUX_s_1_2_2((MUX1HOT_s_1_1_2(1'b1, fsm_output[0])), (MUX1HOT_s_1_1_2(1'b1,
      and_6_nl)), fsm_output[1]);
  assign IsInf_6U_23U_land_lpi_1_dfm_mx1w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm!=10'b0000000000) |
      IsNaN_6U_23U_IsNaN_6U_23U_nand_cse);
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      (chn_a_rsci_d_mxwt[9:0]), IsNaN_6U_23U_land_lpi_1_dfm);
  assign IsNaN_6U_23U_nor_tmp = ~((chn_a_rsci_d_mxwt[9:0]!=10'b0000000000));
  assign IsNaN_6U_23U_land_lpi_1_dfm = ~(IsNaN_6U_23U_nor_tmp | IsNaN_6U_23U_IsNaN_6U_23U_nand_cse);
  assign IsNaN_6U_23U_aelse_not_2_nl = ~ IsNaN_6U_23U_land_lpi_1_dfm;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      (chn_a_rsci_d_mxwt[9:0]), (IsNaN_6U_23U_aelse_not_2_nl));
  assign IsNaN_6U_23U_IsNaN_6U_23U_nand_cse = ~((chn_a_rsci_d_mxwt[15:10]==6'b111111));
  assign or_cse = chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse);
  assign and_4_mdf = chn_a_rsci_bawt & or_cse;
  assign and_dcpl_2 = chn_o_rsci_bawt & reg_chn_o_rsci_ld_core_psct_cse;
  assign or_dcpl_3 = ~((~((~ chn_o_rsci_bawt) & reg_chn_o_rsci_ld_core_psct_cse))
      & chn_a_rsci_bawt);
  assign and_dcpl_7 = (chn_a_rsci_d_mxwt[14:13]==2'b11);
  assign and_dcpl_11 = (chn_a_rsci_d_mxwt[12:10]==3'b111);
  assign or_dcpl_9 = (chn_a_rsci_d_mxwt[15:10]!=6'b111111) | IsNaN_6U_23U_nor_tmp;
  assign and_dcpl_25 = and_dcpl_2 & (~ chn_a_rsci_bawt);
  assign and_46_cse = and_dcpl_11 & or_cse & and_dcpl_7 & (chn_a_rsci_d_mxwt[15])
      & (~ IsNaN_6U_23U_nor_tmp) & chn_a_rsci_bawt & (fsm_output[1]);
  assign and_48_cse = or_dcpl_9 & or_cse & chn_a_rsci_bawt & (fsm_output[1]);
  assign or_tmp_18 = or_cse & chn_a_rsci_bawt & (fsm_output[1]);
  assign chn_a_rsci_ld_core_psct_mx0c0 = and_4_mdf | (fsm_output[0]);
  assign chn_o_rsci_d_9_0_mx0c1 = and_48_cse | (or_dcpl_9 & and_dcpl_2 & chn_a_rsci_bawt);
  assign chn_a_rsci_oswt_unreg = or_tmp_18;
  assign chn_o_rsci_oswt_unreg = and_dcpl_2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_iswt0 <= 1'b0;
      reg_chn_o_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_a_rsci_iswt0 <= ~((~ and_4_mdf) & (fsm_output[1]));
      reg_chn_o_rsci_iswt0_cse <= or_tmp_18;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_a_rsci_ld_core_psct_mx0c0 ) begin
      chn_a_rsci_ld_core_psct <= chn_a_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_10 <= 1'b0;
    end
    else if ( core_wen & (~ (fsm_output[0])) & (~ or_dcpl_3) ) begin
      chn_o_rsci_d_10 <= IsInf_6U_23U_land_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_9_0 <= 10'b0;
    end
    else if ( core_wen & (and_46_cse | (and_dcpl_11 & and_dcpl_7 & (chn_a_rsci_d_mxwt[15])
        & (~ IsNaN_6U_23U_nor_tmp) & chn_o_rsci_bawt & reg_chn_o_rsci_ld_core_psct_cse
        & chn_a_rsci_bawt) | chn_o_rsci_d_9_0_mx0c1) ) begin
      chn_o_rsci_d_9_0 <= MUX_v_10_2_2(({{9{IsInf_6U_23U_land_lpi_1_dfm_mx1w0}},
          IsInf_6U_23U_land_lpi_1_dfm_mx1w0}), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm,
          nand_11_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_22_13 <= 10'b0;
    end
    else if ( core_wen & (and_46_cse | and_48_cse) ) begin
      chn_o_rsci_d_22_13 <= MUX_v_10_2_2(({{9{IsInf_6U_23U_land_lpi_1_dfm_mx1w0}},
          IsInf_6U_23U_land_lpi_1_dfm_mx1w0}), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm,
          nand_10_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_27_23 <= 5'b0;
    end
    else if ( core_wen & (~(or_dcpl_3 | ((~(chn_o_rsci_bawt & reg_chn_o_rsci_ld_core_psct_cse
        & chn_a_rsci_bawt)) & (fsm_output[0])))) ) begin
      chn_o_rsci_d_27_23 <= MUX_v_5_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_mux_5_nl),
          5'b11111, IsNaN_6U_23U_land_lpi_1_dfm);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_30_28 <= 3'b0;
      chn_o_rsci_d_31 <= 1'b0;
    end
    else if ( chn_o_and_4_cse ) begin
      chn_o_rsci_d_30_28 <= (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_nl)
          | ({{2{IsInf_6U_23U_land_lpi_1_dfm_mx1w0}}, IsInf_6U_23U_land_lpi_1_dfm_mx1w0})
          | ({{2{IsNaN_6U_23U_land_lpi_1_dfm}}, IsNaN_6U_23U_land_lpi_1_dfm});
      chn_o_rsci_d_31 <= chn_a_rsci_d_mxwt[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_18 | and_dcpl_25) ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= ~ and_dcpl_25;
    end
  end
  assign nand_11_nl = ~(IsInf_6U_23U_land_lpi_1_dfm_mx1w0 & chn_o_rsci_d_9_0_mx0c1);
  assign nand_10_nl = ~(IsInf_6U_23U_land_lpi_1_dfm_mx1w0 & and_48_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_mux_5_nl = MUX_v_5_2_2((chn_a_rsci_d_mxwt[14:10]),
      5'b11110, IsInf_6U_23U_land_lpi_1_dfm_mx1w0);
  assign nl_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = conv_u2u_2_3({1'b1 , (chn_a_rsci_d_mxwt[15])})
      + 3'b1;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = nl_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl[2:0];
  assign IsZero_6U_23U_aelse_IsZero_6U_23U_or_nl = (chn_a_rsci_d_mxwt[15:0]!=16'b0000000000000000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_nl = MUX_v_3_2_2(3'b000,
      (FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl), (IsZero_6U_23U_aelse_IsZero_6U_23U_or_nl));

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_to_fp32
// ------------------------------------------------------------------


module HLS_fp17_to_fp32 (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_o_rsc_z,
      chn_o_rsc_vz, chn_o_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  output [31:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;


  // Interconnect Declarations
  wire chn_a_rsci_oswt;
  wire chn_a_rsci_oswt_unreg;
  wire chn_o_rsci_oswt;
  wire chn_o_rsci_oswt_unreg;


  // Interconnect Declarations for Component Instantiations 
  FP17_TO_FP32_chn_a_rsci_unreg chn_a_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg),
      .outsig(chn_a_rsci_oswt)
    );
  FP17_TO_FP32_chn_o_rsci_unreg chn_o_rsci_unreg_inst (
      .in_0(chn_o_rsci_oswt_unreg),
      .outsig(chn_o_rsci_oswt)
    );
  HLS_fp17_to_fp32_core HLS_fp17_to_fp32_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_oswt_unreg(chn_a_rsci_oswt_unreg),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_oswt_unreg(chn_o_rsci_oswt_unreg)
    );
endmodule



