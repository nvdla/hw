// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// nvdla_top sv side SC-SV Adapter 
// This is autogenerated code

`ifndef nvdla_top_sv_interface
`define nvdla_top_sv_interface

interface nvdla_top_sv_interface(wire  nvdla_intr);  
endinterface:nvdla_top_sv_interface 

`endif // nvdla_top_sv_interface


