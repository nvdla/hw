`ifndef _MEM_DEFINE_SVH
`define _MEM_DEFINE_SVH

  `define MEM_ADDR_WIDTH    64

  typedef bit[`MEM_ADDR_WIDTH-1:0] addr_t;

`endif
