// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: HLS_fp32_to_fp16.v

module FP32_TO_FP16_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/FP32_TO_FP16_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module FP32_TO_FP16_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v4.v 
module FP32_TO_FP16_mgc_shift_r_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v 
module FP32_TO_FP16_mgc_shift_l_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-159
//  Generated date: Mon Jul  3 21:37:29 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    FP32_TO_FP16_chn_o_rsci_unreg
// ------------------------------------------------------------------


module FP32_TO_FP16_chn_o_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP32_TO_FP16_chn_a_rsci_unreg
// ------------------------------------------------------------------


module FP32_TO_FP16_chn_a_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for HLS_fp32_to_fp16_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : HLS_fp32_to_fp16_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_staller
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_a_rsci_wen_comp, core_wten, chn_o_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_a_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_o_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_a_rsci_wen_comp & chn_o_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_dp
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_biwt, chn_o_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_biwt;
  input chn_o_rsci_bdwt;


  // Interconnect Declarations
  reg chn_o_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_bawt = chn_o_rsci_biwt | chn_o_rsci_bcwt;
  assign chn_o_rsci_wen_comp = (~ chn_o_rsci_oswt) | chn_o_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_o_rsci_bcwt <= ~((~(chn_o_rsci_bcwt | chn_o_rsci_biwt)) | chn_o_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, core_wen, core_wten, chn_o_rsci_iswt0,
      chn_o_rsci_ld_core_psct, chn_o_rsci_biwt, chn_o_rsci_bdwt, chn_o_rsci_ld_core_sct,
      chn_o_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  input chn_o_rsci_ld_core_psct;
  output chn_o_rsci_biwt;
  output chn_o_rsci_bdwt;
  output chn_o_rsci_ld_core_sct;
  input chn_o_rsci_vd;


  // Interconnect Declarations
  wire chn_o_rsci_ogwt;
  wire chn_o_rsci_pdswt0;
  reg chn_o_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_pdswt0 = (~ core_wten) & chn_o_rsci_iswt0;
  assign chn_o_rsci_biwt = chn_o_rsci_ogwt & chn_o_rsci_vd;
  assign chn_o_rsci_ogwt = chn_o_rsci_pdswt0 | chn_o_rsci_icwt;
  assign chn_o_rsci_bdwt = chn_o_rsci_oswt & core_wen;
  assign chn_o_rsci_ld_core_sct = chn_o_rsci_ld_core_psct & chn_o_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_icwt <= 1'b0;
    end
    else begin
      chn_o_rsci_icwt <= ~((~(chn_o_rsci_icwt | chn_o_rsci_pdswt0)) | chn_o_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_dp
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, chn_a_rsci_bawt, chn_a_rsci_wen_comp,
      chn_a_rsci_d_mxwt, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  output [31:0] chn_a_rsci_d_mxwt;
  input chn_a_rsci_biwt;
  input chn_a_rsci_bdwt;
  input [31:0] chn_a_rsci_d;


  // Interconnect Declarations
  reg chn_a_rsci_bcwt;
  reg [31:0] chn_a_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_bawt = chn_a_rsci_biwt | chn_a_rsci_bcwt;
  assign chn_a_rsci_wen_comp = (~ chn_a_rsci_oswt) | chn_a_rsci_bawt;
  assign chn_a_rsci_d_mxwt = MUX_v_32_2_2(chn_a_rsci_d, chn_a_rsci_d_bfwt, chn_a_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_bcwt <= 1'b0;
      chn_a_rsci_d_bfwt <= 32'b0;
    end
    else begin
      chn_a_rsci_bcwt <= ~((~(chn_a_rsci_bcwt | chn_a_rsci_biwt)) | chn_a_rsci_bdwt);
      chn_a_rsci_d_bfwt <= chn_a_rsci_d_mxwt;
    end
  end

  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct,
      core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  input chn_a_rsci_ld_core_psct;
  input core_wten;
  output chn_a_rsci_biwt;
  output chn_a_rsci_bdwt;
  output chn_a_rsci_ld_core_sct;
  input chn_a_rsci_vd;


  // Interconnect Declarations
  wire chn_a_rsci_ogwt;
  wire chn_a_rsci_pdswt0;
  reg chn_a_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_pdswt0 = (~ core_wten) & chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & chn_a_rsci_vd;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | chn_a_rsci_icwt;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & chn_a_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_icwt <= 1'b0;
    end
    else begin
      chn_a_rsci_icwt <= ~((~(chn_a_rsci_icwt | chn_a_rsci_pdswt0)) | chn_a_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_chn_o_rsci
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_chn_o_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_o_rsci_oswt,
      core_wen, core_wten, chn_o_rsci_iswt0, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_ld_core_psct, chn_o_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [15:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_ld_core_psct;
  input [15:0] chn_o_rsci_d;


  // Interconnect Declarations
  wire chn_o_rsci_biwt;
  wire chn_o_rsci_bdwt;
  wire chn_o_rsci_ld_core_sct;
  wire chn_o_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  FP32_TO_FP16_mgc_out_stdreg_wait_v1 #(.rscid(32'sd2),
  .width(32'sd16)) chn_o_rsci (
      .ld(chn_o_rsci_ld_core_sct),
      .vd(chn_o_rsci_vd),
      .d(chn_o_rsci_d),
      .lz(chn_o_rsc_lz),
      .vz(chn_o_rsc_vz),
      .z(chn_o_rsc_z)
    );
  HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_ctrl HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_ld_core_psct(chn_o_rsci_ld_core_psct),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt),
      .chn_o_rsci_ld_core_sct(chn_o_rsci_ld_core_sct),
      .chn_o_rsci_vd(chn_o_rsci_vd)
    );
  HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_dp HLS_fp32_to_fp16_core_chn_o_rsci_chn_o_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core_chn_a_rsci
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core_chn_a_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_a_rsci_oswt,
      core_wen, chn_a_rsci_iswt0, chn_a_rsci_bawt, chn_a_rsci_wen_comp, chn_a_rsci_ld_core_psct,
      chn_a_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  input chn_a_rsci_ld_core_psct;
  output [31:0] chn_a_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_a_rsci_biwt;
  wire chn_a_rsci_bdwt;
  wire chn_a_rsci_ld_core_sct;
  wire chn_a_rsci_vd;
  wire [31:0] chn_a_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP32_TO_FP16_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd32)) chn_a_rsci (
      .ld(chn_a_rsci_ld_core_sct),
      .vd(chn_a_rsci_vd),
      .d(chn_a_rsci_d),
      .lz(chn_a_rsc_lz),
      .vz(chn_a_rsc_vz),
      .z(chn_a_rsc_z)
    );
  HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_ctrl HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_ld_core_sct(chn_a_rsci_ld_core_sct),
      .chn_a_rsci_vd(chn_a_rsci_vd)
    );
  HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_dp HLS_fp32_to_fp16_core_chn_a_rsci_chn_a_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_d(chn_a_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16_core
// ------------------------------------------------------------------


module HLS_fp32_to_fp16_core (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_o_rsc_z,
      chn_o_rsc_vz, chn_o_rsc_lz, chn_a_rsci_oswt, chn_a_rsci_oswt_unreg, chn_o_rsci_oswt,
      chn_o_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  output [15:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_a_rsci_oswt;
  output chn_a_rsci_oswt_unreg;
  input chn_o_rsci_oswt;
  output chn_o_rsci_oswt_unreg;


  // Interconnect Declarations
  wire core_wen;
  reg chn_a_rsci_iswt0;
  wire chn_a_rsci_bawt;
  wire chn_a_rsci_wen_comp;
  reg chn_a_rsci_ld_core_psct;
  wire [31:0] chn_a_rsci_d_mxwt;
  wire core_wten;
  reg chn_o_rsci_iswt0;
  wire chn_o_rsci_bawt;
  wire chn_o_rsci_wen_comp;
  reg chn_o_rsci_d_15;
  reg [9:0] chn_o_rsci_d_9_0;
  reg chn_o_rsci_d_14;
  reg [3:0] chn_o_rsci_d_13_10;
  wire [1:0] fsm_output;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nand_tmp;
  wire IsNaN_8U_23U_nor_tmp;
  wire or_tmp_2;
  wire mux_tmp;
  wire mux_tmp_1;
  wire and_tmp;
  wire or_tmp_7;
  wire or_tmp_9;
  wire or_tmp_25;
  wire or_tmp_26;
  wire mux_tmp_16;
  wire mux_tmp_19;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_28;
  wire or_dcpl_11;
  wire or_tmp_53;
  reg FpMantRNE_24U_11U_else_and_svs;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2;
  reg FpMantRNE_24U_11U_else_carry_sva_2;
  reg FpMantRNE_24U_11U_else_and_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5;
  reg IsNaN_8U_23U_land_lpi_1_dfm_2;
  reg [10:0] FpMantDecShiftRight_23U_8U_10U_i_mant_s_slc_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_23_13_itm_2;
  reg FpMantDecShiftRight_23U_8U_10U_carry_and_itm_2;
  reg IsNaN_8U_23U_nor_itm_2;
  reg IsNaN_8U_23U_IsNaN_8U_23U_nand_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_4;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_4;
  reg FpMantRNE_24U_11U_else_and_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_31_1;
  reg [27:0] FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_31_1;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_9_0_1;
  wire main_stage_en_1;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp;
  wire FpMantRNE_24U_11U_else_carry_sva_mx0w0;
  wire [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4;
  wire [5:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4;
  wire chn_o_and_cse;
  wire or_7_cse;
  wire nor_15_cse;
  wire and_72_cse;
  reg reg_chn_o_rsci_ld_core_psct_cse;
  wire and_74_cse;
  wire nor_2_cse;
  wire and_37_cse;
  wire and_43_rgt;
  wire and_49_rgt;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  wire FpMantDecShiftRight_23U_8U_10U_stick_mask_and_tmp;
  wire [22:0] z_out;
  wire [23:0] nl_z_out;
  wire HLS_fp32_to_fp16_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_sig_mx0;
  wire chn_a_rsci_ld_core_psct_mx0c0;
  wire chn_o_rsci_d_9_0_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire FpMantRNE_24U_11U_else_and_svs_mx0w0;
  wire main_stage_v_2_mx0c1;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_sva;
  wire [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva;
  wire FpMantDecShiftRight_23U_8U_10U_i_mant_s_and_cse;
  wire Fp32ToFp16_and_1_cse;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_if_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_or_cse;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1;

  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] shift_0_prb;
  wire[0:0] and_11;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_2_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] or_2_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] and_76_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] or_12_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_15_nl;
  wire[0:0] nor_25_nl;
  wire[0:0] nor_4_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] nor_5_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] nor_34_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_19_nl;
  wire[0:0] and_73_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] nor_17_nl;
  wire[0:0] nor_18_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] and_70_nl;
  wire[0:0] and_19_nl;
  wire[8:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  wire[9:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  wire[8:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  wire[8:0] FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  wire[9:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] and_75_nl;
  wire[22:0] FpMantRNE_24U_11U_else_mux_4_nl;
  wire[0:0] FpMantRNE_24U_11U_else_FpMantRNE_24U_11U_else_or_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  assign nl_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = {1'b1 , (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[22:0])};
  wire [3:0] nl_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  assign nl_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[23]))};
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva
      + 5'b11111;
  wire [15:0] nl_HLS_fp32_to_fp16_core_chn_o_rsci_inst_chn_o_rsci_d;
  assign nl_HLS_fp32_to_fp16_core_chn_o_rsci_inst_chn_o_rsci_d = {chn_o_rsci_d_15
      , chn_o_rsci_d_14 , chn_o_rsci_d_13_10 , chn_o_rsci_d_9_0};
  FP32_TO_FP16_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg (
      .a(nl_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a[23:0]),
      .s(nl_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
    );
  FP32_TO_FP16_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg (
      .a(1'b1),
      .s(nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_sva)
    );
  FP32_TO_FP16_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_sva)
    );
  HLS_fp32_to_fp16_core_chn_a_rsci HLS_fp32_to_fp16_core_chn_a_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  HLS_fp32_to_fp16_core_chn_o_rsci HLS_fp32_to_fp16_core_chn_o_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_ld_core_psct(reg_chn_o_rsci_ld_core_psct_cse),
      .chn_o_rsci_d(nl_HLS_fp32_to_fp16_core_chn_o_rsci_inst_chn_o_rsci_d[15:0])
    );
  HLS_fp32_to_fp16_core_staller HLS_fp32_to_fp16_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp)
    );
  HLS_fp32_to_fp16_core_core_fsm HLS_fp32_to_fp16_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign iMantWidth_oMantWidth_prb = HLS_fp32_to_fp16_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_sig_mx0;
  // assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
  // PSL HLS_fp32_to_fp16_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb = HLS_fp32_to_fp16_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_sig_mx0;
  // assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
  // PSL HLS_fp32_to_fp16_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign and_11 = and_37_cse & FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3);
  assign shift_0_prb = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2)
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[23])}) + 5'b1)), and_11);
  // assert(shift > 0) - ../include/nvdla_float.h: line 286
  // PSL HLS_fp32_to_fp16_core_nvdla_float_h_ln286_assert_shift_gt_0 : assert { shift_0_prb } @rose(nvdla_core_clk);
  assign chn_o_and_cse = core_wen & (~(and_dcpl_8 | (~ main_stage_v_2)));
  assign or_7_cse = (~ reg_chn_o_rsci_ld_core_psct_cse) | chn_o_rsci_bawt;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse = core_wen & (~ and_dcpl_8) &
      mux_tmp;
  assign and_37_cse = or_7_cse & main_stage_v_1;
  assign nor_21_nl = ~((~ or_tmp_9) | (~ main_stage_v_1) | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3);
  assign nor_34_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4
      | (~ main_stage_v_2) | IsNaN_8U_23U_land_lpi_1_dfm_2 | FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_4
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_4
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4);
  assign mux_14_nl = MUX_s_1_2_2((nor_34_nl), (nor_21_nl), or_7_cse);
  assign FpMantDecShiftRight_23U_8U_10U_i_mant_s_and_cse = core_wen & (~ and_dcpl_8)
      & (mux_14_nl);
  assign Fp32ToFp16_and_1_cse = core_wen & (~ and_dcpl_8) & mux_tmp_19;
  assign nor_15_cse = ~(IsNaN_8U_23U_IsNaN_8U_23U_nand_itm_2 | IsNaN_8U_23U_nor_itm_2);
  assign and_72_cse = (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4==5'b11111) & FpMantRNE_24U_11U_else_and_svs_2;
  assign and_74_cse = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4
      & FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4;
  assign and_43_rgt = or_7_cse & or_tmp_9;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_if_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_or_cse
      = (or_7_cse & FpMantRNE_24U_11U_else_and_svs_2) | and_dcpl_28;
  assign and_49_rgt = or_dcpl_11 & or_7_cse;
  assign and_19_nl = main_stage_en_1 & (fsm_output[1]);
  assign HLS_fp32_to_fp16_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_sig_mx0
      = MUX_s_1_2_2((MUX1HOT_s_1_1_2(1'b1, fsm_output[0])), (MUX1HOT_s_1_1_2(1'b1,
      and_19_nl)), fsm_output[1]);
  assign FpMantRNE_24U_11U_else_and_svs_mx0w0 = FpMantRNE_24U_11U_else_carry_sva_mx0w0
      & (chn_a_rsci_d_mxwt[22:13]==10'b1111111111);
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1 , (~ (chn_a_rsci_d_mxwt[30:23]))})
      + 9'b1110001;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1 = readslicef_9_1_8((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_7_8(chn_a_rsci_d_mxwt[30:24])
      + 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 = readslicef_8_1_7((FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl = conv_u2s_8_9(chn_a_rsci_d_mxwt[30:23])
      + 9'b101110001;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1 = readslicef_9_1_8((FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl));
  assign FpMantRNE_24U_11U_else_carry_sva_mx0w0 = (chn_a_rsci_d_mxwt[12]) & ((chn_a_rsci_d_mxwt[0])
      | (chn_a_rsci_d_mxwt[1]) | (chn_a_rsci_d_mxwt[2]) | (chn_a_rsci_d_mxwt[3])
      | (chn_a_rsci_d_mxwt[4]) | (chn_a_rsci_d_mxwt[5]) | (chn_a_rsci_d_mxwt[6])
      | (chn_a_rsci_d_mxwt[7]) | (chn_a_rsci_d_mxwt[8]) | (chn_a_rsci_d_mxwt[9])
      | (chn_a_rsci_d_mxwt[10]) | (chn_a_rsci_d_mxwt[11]) | (chn_a_rsci_d_mxwt[13]));
  assign IsNaN_8U_23U_nor_tmp = ~((chn_a_rsci_d_mxwt[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_IsNaN_8U_23U_nand_tmp = ~((chn_a_rsci_d_mxwt[30:23]==8'b11111111));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = FpMantDecShiftRight_23U_8U_10U_i_mant_s_slc_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_23_13_itm_2
      + conv_u2u_1_11(FpMantDecShiftRight_23U_8U_10U_carry_and_itm_2);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc =
      ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp | FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4);
  assign main_stage_en_1 = chn_a_rsci_bawt & or_7_cse;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4 = ({(~ (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[27]))
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[26:23])}) + 5'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4 = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4[4:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva = (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[22:0])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0]);
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva = (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[22:0])
      & z_out;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva = (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[22:0])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_sva[22:0]);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[23]))}) + 5'b1101;
  assign FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva = nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva[4:0];
  assign or_tmp_2 = chn_o_rsci_bawt | (~(reg_chn_o_rsci_ld_core_psct_cse & main_stage_v_1));
  assign nor_2_cse = ~(chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign mux_tmp = MUX_s_1_2_2(chn_a_rsci_bawt, main_stage_v_1, nor_2_cse);
  assign mux_tmp_1 = MUX_s_1_2_2((~ or_tmp_2), mux_tmp, FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1);
  assign nor_28_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ chn_a_rsci_bawt));
  assign mux_3_nl = MUX_s_1_2_2((nor_28_nl), chn_a_rsci_bawt, chn_o_rsci_bawt);
  assign and_tmp = FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1 & (mux_3_nl);
  assign or_tmp_7 = IsNaN_8U_23U_IsNaN_8U_23U_nand_tmp | IsNaN_8U_23U_nor_tmp;
  assign or_tmp_9 = IsNaN_8U_23U_nor_itm_2 | IsNaN_8U_23U_IsNaN_8U_23U_nand_itm_2;
  assign or_tmp_25 = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4
      & main_stage_v_2 & (~ chn_o_rsci_bawt) & reg_chn_o_rsci_ld_core_psct_cse);
  assign or_tmp_26 = nor_2_cse | main_stage_v_1;
  assign and_75_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4
      & main_stage_v_2;
  assign mux_15_nl = MUX_s_1_2_2(and_37_cse, or_tmp_26, and_75_nl);
  assign mux_tmp_16 = MUX_s_1_2_2((~ or_tmp_25), (mux_15_nl), FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3);
  assign mux_tmp_19 = MUX_s_1_2_2(and_37_cse, or_tmp_26, main_stage_v_2);
  assign and_dcpl_6 = reg_chn_o_rsci_ld_core_psct_cse & chn_o_rsci_bawt;
  assign and_dcpl_8 = reg_chn_o_rsci_ld_core_psct_cse & (~ chn_o_rsci_bawt);
  assign and_dcpl_14 = or_7_cse & main_stage_v_2;
  assign and_dcpl_15 = and_dcpl_6 & (~ main_stage_v_2);
  assign and_dcpl_28 = or_7_cse & (~ FpMantRNE_24U_11U_else_and_svs_2);
  assign or_dcpl_11 = (~ FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1) | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1);
  assign or_tmp_53 = or_7_cse & chn_a_rsci_bawt & (fsm_output[1]);
  assign chn_a_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign chn_o_rsci_d_9_0_mx0c1 = or_7_cse & main_stage_v_2 & (~ IsNaN_8U_23U_land_lpi_1_dfm_2);
  assign main_stage_v_1_mx0c1 = or_7_cse & main_stage_v_1 & (~ chn_a_rsci_bawt);
  assign main_stage_v_2_mx0c1 = or_7_cse & (~ main_stage_v_1) & main_stage_v_2;
  assign chn_a_rsci_oswt_unreg = or_tmp_53;
  assign chn_o_rsci_oswt_unreg = and_dcpl_6;
  assign FpMantDecShiftRight_23U_8U_10U_stick_mask_and_tmp = (fsm_output[1]) & (~
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_iswt0 <= 1'b0;
      chn_o_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_a_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_o_rsci_iswt0 <= and_dcpl_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_a_rsci_ld_core_psct_mx0c0 ) begin
      chn_a_rsci_ld_core_psct <= chn_a_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_13_10 <= 4'b0;
      chn_o_rsci_d_14 <= 1'b0;
      chn_o_rsci_d_15 <= 1'b0;
    end
    else if ( chn_o_and_cse ) begin
      chn_o_rsci_d_13_10 <= MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl),
          4'b1111, IsNaN_8U_23U_land_lpi_1_dfm_2);
      chn_o_rsci_d_14 <= (~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_4_1
          & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc))
          | FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5)) | and_74_cse)) |
          IsNaN_8U_23U_land_lpi_1_dfm_2;
      chn_o_rsci_d_15 <= FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_31_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_9_0 <= 10'b0;
    end
    else if ( core_wen & ((or_7_cse & main_stage_v_2 & IsNaN_8U_23U_land_lpi_1_dfm_2)
        | chn_o_rsci_d_9_0_mx0c1) ) begin
      chn_o_rsci_d_9_0 <= MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_9_0_1,
          (FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl),
          chn_o_rsci_d_9_0_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_14 | and_dcpl_15) ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= ~ and_dcpl_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_53 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_4_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 <= nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2[2:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1 <= 28'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_7_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1 <= chn_a_rsci_d_mxwt[27:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_9_nl) ) begin
      FpMantRNE_24U_11U_else_and_svs_st_2 <= FpMantRNE_24U_11U_else_and_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_11_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_12_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_31_1 <= 1'b0;
      IsNaN_8U_23U_nor_itm_2 <= 1'b0;
      IsNaN_8U_23U_IsNaN_8U_23U_nand_itm_2 <= 1'b0;
    end
    else if ( FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_31_1 <= chn_a_rsci_d_mxwt[31];
      IsNaN_8U_23U_nor_itm_2 <= IsNaN_8U_23U_nor_tmp;
      IsNaN_8U_23U_IsNaN_8U_23U_nand_itm_2 <= IsNaN_8U_23U_IsNaN_8U_23U_nand_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_37_cse | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_i_mant_s_slc_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_23_13_itm_2
          <= 11'b0;
      FpMantDecShiftRight_23U_8U_10U_carry_and_itm_2 <= 1'b0;
    end
    else if ( FpMantDecShiftRight_23U_8U_10U_i_mant_s_and_cse ) begin
      FpMantDecShiftRight_23U_8U_10U_i_mant_s_slc_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_23_13_itm_2
          <= FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13];
      FpMantDecShiftRight_23U_8U_10U_carry_and_itm_2 <= ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva!=23'b00000000000000000000000)
          | (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva!=23'b00000000000000000000000)
          | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva!=23'b00000000000000000000000)
          | (FpMantDecShiftRight_23U_8U_10U_least_mask_sva[23]));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_18_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_4
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & mux_tmp_16 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_4
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_31_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_2 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4
          <= 1'b0;
    end
    else if ( Fp32ToFp16_and_1_cse ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_31_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_31_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3;
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4==5'b11111)
          & FpMantRNE_24U_11U_else_and_svs_2 & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3
          & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3)))
          & FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3);
      IsNaN_8U_23U_land_lpi_1_dfm_2 <= nor_15_cse;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3;
      FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_4
          <= FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_9_0_1 <= 10'b0;
    end
    else if ( core_wen & ((or_7_cse & nor_15_cse) | and_43_rgt) & (mux_21_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_9_0_1 <= MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[9:0]),
          (z_out[9:0]), and_43_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_4_1 <= 1'b0;
    end
    else if ( core_wen & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_if_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_or_cse
        & mux_tmp_19 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_4_1 <= MUX_s_1_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4[4]),
          (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[27])), and_dcpl_28);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_3_0_1 <= 4'b0;
    end
    else if ( core_wen & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_if_FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_or_cse
        & (mux_22_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_3_0_1 <= MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_4[3:0]),
          (FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[26:23]), and_dcpl_28);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_7_cse & FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1
        & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1) & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1)
        | and_49_rgt) & mux_tmp ) begin
      FpMantRNE_24U_11U_else_and_svs_2 <= MUX_s_1_2_2(FpMantRNE_24U_11U_else_and_svs_mx0w0,
          FpMantRNE_24U_11U_else_and_svs, and_49_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_8) & (mux_23_nl) ) begin
      FpMantRNE_24U_11U_else_carry_sva_2 <= FpMantRNE_24U_11U_else_carry_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_8 | (~ chn_a_rsci_bawt) | or_dcpl_11 | (fsm_output[0])))
        ) begin
      FpMantRNE_24U_11U_else_and_svs <= FpMantRNE_24U_11U_else_and_svs_mx0w0;
    end
  end
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl =
      MUX1HOT_v_4_3_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10])}),
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_8_3_0_1, 4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_nl) , FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_2_nl = ~ and_74_cse;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_2_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[9:0]),
      FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_2_9_0_1, FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl),
      10'b1111111111, FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl), 10'b1111111111,
      and_74_cse));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 
      = (~ (chn_a_rsci_d_mxwt[26:24])) + 3'b1;
  assign or_2_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1 | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
  assign mux_2_nl = MUX_s_1_2_2(mux_tmp_1, (~ or_tmp_2), or_2_nl);
  assign nor_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1 | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1
      | (~ and_tmp));
  assign nor_31_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3));
  assign mux_4_nl = MUX_s_1_2_2((nor_nl), (mux_2_nl), nor_31_nl);
  assign and_76_nl = chn_a_rsci_bawt & (~(or_tmp_7 & (FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1))));
  assign nor_27_nl = ~(FpMantRNE_24U_11U_else_and_svs_2 | (~ main_stage_v_1));
  assign or_12_nl = (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3)))
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3)
      | FpMantRNE_24U_11U_else_and_svs_st_2;
  assign mux_5_nl = MUX_s_1_2_2((nor_27_nl), main_stage_v_1, or_12_nl);
  assign nor_26_nl = ~((~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
      | (~ (mux_5_nl)));
  assign mux_6_nl = MUX_s_1_2_2(main_stage_v_1, (nor_26_nl), or_tmp_9);
  assign mux_7_nl = MUX_s_1_2_2((mux_6_nl), (and_76_nl), or_7_cse);
  assign or_15_nl = (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1) | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
  assign mux_8_nl = MUX_s_1_2_2(mux_tmp_1, (~ or_tmp_2), or_15_nl);
  assign nor_25_nl = ~((~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1) |
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~ and_tmp));
  assign nor_4_nl = ~((~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3));
  assign mux_9_nl = MUX_s_1_2_2((nor_25_nl), (mux_8_nl), nor_4_nl);
  assign mux_10_nl = MUX_s_1_2_2(mux_tmp_1, (~ or_tmp_2), FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1);
  assign nor_24_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~ and_tmp));
  assign nor_5_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3));
  assign mux_11_nl = MUX_s_1_2_2((nor_24_nl), (mux_10_nl), nor_5_nl);
  assign mux_12_nl = MUX_s_1_2_2(and_tmp, mux_tmp_1, FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3);
  assign nor_20_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3
      | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3
      & and_37_cse)));
  assign mux_17_nl = MUX_s_1_2_2(mux_tmp_16, (~ or_tmp_25), FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3);
  assign mux_18_nl = MUX_s_1_2_2((mux_17_nl), (nor_20_nl), FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_4);
  assign nor_19_nl = ~(and_72_cse | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3
      | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3
      & main_stage_v_1)));
  assign mux_20_nl = MUX_s_1_2_2(main_stage_v_1, (nor_19_nl), or_tmp_9);
  assign and_73_nl = ((~(and_74_cse | FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4)))
      | IsNaN_8U_23U_land_lpi_1_dfm_2) & main_stage_v_2;
  assign mux_21_nl = MUX_s_1_2_2((and_73_nl), (mux_20_nl), or_7_cse);
  assign nor_17_nl = ~(and_72_cse | (~(or_tmp_9 & main_stage_v_1 & FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3)));
  assign nor_18_nl = ~((~ main_stage_v_2) | IsNaN_8U_23U_land_lpi_1_dfm_2 | FpWidthDec_8U_23U_5U_10U_1U_1U_is_inf_lpi_1_dfm_5
      | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_4)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_4);
  assign mux_22_nl = MUX_s_1_2_2((nor_18_nl), (nor_17_nl), or_7_cse);
  assign nor_16_nl = ~((~ or_tmp_7) | (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1
      & chn_a_rsci_bawt)));
  assign and_70_nl = or_tmp_9 & main_stage_v_1 & FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_3
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_3)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_3
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_3)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_3;
  assign mux_23_nl = MUX_s_1_2_2((and_70_nl), (nor_16_nl), or_7_cse);
  assign FpMantRNE_24U_11U_else_mux_4_nl = MUX_v_23_2_2((signext_23_10(FpWidthDec_8U_23U_5U_10U_1U_1U_bits_sva_1_27_0_1[22:13])),
      (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0]), FpMantDecShiftRight_23U_8U_10U_stick_mask_and_tmp);
  assign FpMantRNE_24U_11U_else_FpMantRNE_24U_11U_else_or_2_nl = FpMantRNE_24U_11U_else_carry_sva_2
      | FpMantDecShiftRight_23U_8U_10U_stick_mask_and_tmp;
  assign nl_z_out = (FpMantRNE_24U_11U_else_mux_4_nl) + conv_s2u_2_23({FpMantDecShiftRight_23U_8U_10U_stick_mask_and_tmp
      , (FpMantRNE_24U_11U_else_FpMantRNE_24U_11U_else_or_2_nl)});
  assign z_out = nl_z_out[22:0];

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function [22:0] signext_23_10;
    input [9:0] vector;
  begin
    signext_23_10= {{13{vector[9]}}, vector};
  end
  endfunction


  function  [22:0] conv_s2u_2_23 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_23 = {{21{vector[1]}}, vector};
  end
  endfunction


  function  [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function  [10:0] conv_u2u_1_11 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function  [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp32_to_fp16
// ------------------------------------------------------------------


module HLS_fp32_to_fp16 (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_o_rsc_z,
      chn_o_rsc_vz, chn_o_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [31:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  output [15:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;


  // Interconnect Declarations
  wire chn_a_rsci_oswt;
  wire chn_a_rsci_oswt_unreg;
  wire chn_o_rsci_oswt;
  wire chn_o_rsci_oswt_unreg;


  // Interconnect Declarations for Component Instantiations 
  FP32_TO_FP16_chn_a_rsci_unreg chn_a_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg),
      .outsig(chn_a_rsci_oswt)
    );
  FP32_TO_FP16_chn_o_rsci_unreg chn_o_rsci_unreg_inst (
      .in_0(chn_o_rsci_oswt_unreg),
      .outsig(chn_o_rsci_oswt)
    );
  HLS_fp32_to_fp16_core HLS_fp32_to_fp16_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_oswt_unreg(chn_a_rsci_oswt_unreg),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_oswt_unreg(chn_o_rsci_oswt_unreg)
    );
endmodule



