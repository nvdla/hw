`ifndef _CC_DEFINES_SV_
`define _CC_DEFINES_SV_

//`define CC_MAC2ACCU_DATA_WIDTH   176  
//`define CC_MAC2ACCU_DATA_LENGTH  16
//`define CC_MAC2ACCU_MASK_WIDTH   16
//`define CC_SC2MAC_DATA_WIDTH     8
//`define CC_SC2MAC_DATA_LENGTH    128
//`define CC_SC2MAC_MASK_WIDTH     128
`define CC_PD_WIDTH              9
`define CC_SEL_WIDTH             16

`endif // _CC_DEFINES_SV_
