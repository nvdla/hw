// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_NVDLA_CSC_WL_dec.v

module NV_NVDLA_CSC_WL_dec (
   nvdla_core_clk
  ,nvdla_core_rstn
  ,input_data
  ,input_mask
  ,input_mask_en
  ,input_pipe_valid
  ,input_sel
  ,is_fp16
  ,is_int8
  ,output_data0
  ,output_data1
  ,output_data10
  ,output_data100
  ,output_data101
  ,output_data102
  ,output_data103
  ,output_data104
  ,output_data105
  ,output_data106
  ,output_data107
  ,output_data108
  ,output_data109
  ,output_data11
  ,output_data110
  ,output_data111
  ,output_data112
  ,output_data113
  ,output_data114
  ,output_data115
  ,output_data116
  ,output_data117
  ,output_data118
  ,output_data119
  ,output_data12
  ,output_data120
  ,output_data121
  ,output_data122
  ,output_data123
  ,output_data124
  ,output_data125
  ,output_data126
  ,output_data127
  ,output_data13
  ,output_data14
  ,output_data15
  ,output_data16
  ,output_data17
  ,output_data18
  ,output_data19
  ,output_data2
  ,output_data20
  ,output_data21
  ,output_data22
  ,output_data23
  ,output_data24
  ,output_data25
  ,output_data26
  ,output_data27
  ,output_data28
  ,output_data29
  ,output_data3
  ,output_data30
  ,output_data31
  ,output_data32
  ,output_data33
  ,output_data34
  ,output_data35
  ,output_data36
  ,output_data37
  ,output_data38
  ,output_data39
  ,output_data4
  ,output_data40
  ,output_data41
  ,output_data42
  ,output_data43
  ,output_data44
  ,output_data45
  ,output_data46
  ,output_data47
  ,output_data48
  ,output_data49
  ,output_data5
  ,output_data50
  ,output_data51
  ,output_data52
  ,output_data53
  ,output_data54
  ,output_data55
  ,output_data56
  ,output_data57
  ,output_data58
  ,output_data59
  ,output_data6
  ,output_data60
  ,output_data61
  ,output_data62
  ,output_data63
  ,output_data64
  ,output_data65
  ,output_data66
  ,output_data67
  ,output_data68
  ,output_data69
  ,output_data7
  ,output_data70
  ,output_data71
  ,output_data72
  ,output_data73
  ,output_data74
  ,output_data75
  ,output_data76
  ,output_data77
  ,output_data78
  ,output_data79
  ,output_data8
  ,output_data80
  ,output_data81
  ,output_data82
  ,output_data83
  ,output_data84
  ,output_data85
  ,output_data86
  ,output_data87
  ,output_data88
  ,output_data89
  ,output_data9
  ,output_data90
  ,output_data91
  ,output_data92
  ,output_data93
  ,output_data94
  ,output_data95
  ,output_data96
  ,output_data97
  ,output_data98
  ,output_data99
  ,output_mask
  ,output_pvld
  ,output_sel
  );


input           nvdla_core_clk;
input           nvdla_core_rstn;
input  [1023:0] input_data;
input   [127:0] input_mask;
input     [9:0] input_mask_en;
input           input_pipe_valid;
input    [15:0] input_sel;
input           is_fp16;
input           is_int8;
output    [7:0] output_data0;
output    [7:0] output_data1;
output    [7:0] output_data10;
output    [7:0] output_data100;
output    [7:0] output_data101;
output    [7:0] output_data102;
output    [7:0] output_data103;
output    [7:0] output_data104;
output    [7:0] output_data105;
output    [7:0] output_data106;
output    [7:0] output_data107;
output    [7:0] output_data108;
output    [7:0] output_data109;
output    [7:0] output_data11;
output    [7:0] output_data110;
output    [7:0] output_data111;
output    [7:0] output_data112;
output    [7:0] output_data113;
output    [7:0] output_data114;
output    [7:0] output_data115;
output    [7:0] output_data116;
output    [7:0] output_data117;
output    [7:0] output_data118;
output    [7:0] output_data119;
output    [7:0] output_data12;
output    [7:0] output_data120;
output    [7:0] output_data121;
output    [7:0] output_data122;
output    [7:0] output_data123;
output    [7:0] output_data124;
output    [7:0] output_data125;
output    [7:0] output_data126;
output    [7:0] output_data127;
output    [7:0] output_data13;
output    [7:0] output_data14;
output    [7:0] output_data15;
output    [7:0] output_data16;
output    [7:0] output_data17;
output    [7:0] output_data18;
output    [7:0] output_data19;
output    [7:0] output_data2;
output    [7:0] output_data20;
output    [7:0] output_data21;
output    [7:0] output_data22;
output    [7:0] output_data23;
output    [7:0] output_data24;
output    [7:0] output_data25;
output    [7:0] output_data26;
output    [7:0] output_data27;
output    [7:0] output_data28;
output    [7:0] output_data29;
output    [7:0] output_data3;
output    [7:0] output_data30;
output    [7:0] output_data31;
output    [7:0] output_data32;
output    [7:0] output_data33;
output    [7:0] output_data34;
output    [7:0] output_data35;
output    [7:0] output_data36;
output    [7:0] output_data37;
output    [7:0] output_data38;
output    [7:0] output_data39;
output    [7:0] output_data4;
output    [7:0] output_data40;
output    [7:0] output_data41;
output    [7:0] output_data42;
output    [7:0] output_data43;
output    [7:0] output_data44;
output    [7:0] output_data45;
output    [7:0] output_data46;
output    [7:0] output_data47;
output    [7:0] output_data48;
output    [7:0] output_data49;
output    [7:0] output_data5;
output    [7:0] output_data50;
output    [7:0] output_data51;
output    [7:0] output_data52;
output    [7:0] output_data53;
output    [7:0] output_data54;
output    [7:0] output_data55;
output    [7:0] output_data56;
output    [7:0] output_data57;
output    [7:0] output_data58;
output    [7:0] output_data59;
output    [7:0] output_data6;
output    [7:0] output_data60;
output    [7:0] output_data61;
output    [7:0] output_data62;
output    [7:0] output_data63;
output    [7:0] output_data64;
output    [7:0] output_data65;
output    [7:0] output_data66;
output    [7:0] output_data67;
output    [7:0] output_data68;
output    [7:0] output_data69;
output    [7:0] output_data7;
output    [7:0] output_data70;
output    [7:0] output_data71;
output    [7:0] output_data72;
output    [7:0] output_data73;
output    [7:0] output_data74;
output    [7:0] output_data75;
output    [7:0] output_data76;
output    [7:0] output_data77;
output    [7:0] output_data78;
output    [7:0] output_data79;
output    [7:0] output_data8;
output    [7:0] output_data80;
output    [7:0] output_data81;
output    [7:0] output_data82;
output    [7:0] output_data83;
output    [7:0] output_data84;
output    [7:0] output_data85;
output    [7:0] output_data86;
output    [7:0] output_data87;
output    [7:0] output_data88;
output    [7:0] output_data89;
output    [7:0] output_data9;
output    [7:0] output_data90;
output    [7:0] output_data91;
output    [7:0] output_data92;
output    [7:0] output_data93;
output    [7:0] output_data94;
output    [7:0] output_data95;
output    [7:0] output_data96;
output    [7:0] output_data97;
output    [7:0] output_data98;
output    [7:0] output_data99;
output  [127:0] output_mask;
output          output_pvld;
output   [15:0] output_sel;
wire    [127:0] input_mask_gated;
reg    [1023:0] data_d1;
reg     [127:0] mask_d1;
reg     [127:0] mask_d2_fp16_w;
reg     [127:0] mask_d2_int16_w;
reg     [127:0] mask_d2_int8_w;
reg     [127:0] mask_d2_w;
reg     [127:0] mask_d3;
reg      [15:0] sel_d1;
reg      [15:0] sel_d2;
reg      [15:0] sel_d3;
reg             valid_d1;
reg             valid_d2;
reg             valid_d3;
reg       [7:0] vec_data_000;
reg       [7:0] vec_data_000_d2;
reg       [7:0] vec_data_000_d3;
reg       [7:0] vec_data_001;
reg       [7:0] vec_data_001_d2;
reg       [7:0] vec_data_001_d3;
reg       [7:0] vec_data_002;
reg       [7:0] vec_data_002_d2;
reg       [7:0] vec_data_002_d3;
reg       [7:0] vec_data_003;
reg       [7:0] vec_data_003_d2;
reg       [7:0] vec_data_003_d3;
reg       [7:0] vec_data_004;
reg       [7:0] vec_data_004_d2;
reg       [7:0] vec_data_004_d3;
reg       [7:0] vec_data_005;
reg       [7:0] vec_data_005_d2;
reg       [7:0] vec_data_005_d3;
reg       [7:0] vec_data_006;
reg       [7:0] vec_data_006_d2;
reg       [7:0] vec_data_006_d3;
reg       [7:0] vec_data_007;
reg       [7:0] vec_data_007_d2;
reg       [7:0] vec_data_007_d3;
reg       [7:0] vec_data_008;
reg       [7:0] vec_data_008_d2;
reg       [7:0] vec_data_008_d3;
reg       [7:0] vec_data_009;
reg       [7:0] vec_data_009_d2;
reg       [7:0] vec_data_009_d3;
reg       [7:0] vec_data_010;
reg       [7:0] vec_data_010_d2;
reg       [7:0] vec_data_010_d3;
reg       [7:0] vec_data_011;
reg       [7:0] vec_data_011_d2;
reg       [7:0] vec_data_011_d3;
reg       [7:0] vec_data_012;
reg       [7:0] vec_data_012_d2;
reg       [7:0] vec_data_012_d3;
reg       [7:0] vec_data_013;
reg       [7:0] vec_data_013_d2;
reg       [7:0] vec_data_013_d3;
reg       [7:0] vec_data_014;
reg       [7:0] vec_data_014_d2;
reg       [7:0] vec_data_014_d3;
reg       [7:0] vec_data_015;
reg       [7:0] vec_data_015_d2;
reg       [7:0] vec_data_015_d3;
reg       [7:0] vec_data_016;
reg       [7:0] vec_data_016_d2;
reg       [7:0] vec_data_016_d3;
reg       [7:0] vec_data_017;
reg       [7:0] vec_data_017_d2;
reg       [7:0] vec_data_017_d3;
reg       [7:0] vec_data_018;
reg       [7:0] vec_data_018_d2;
reg       [7:0] vec_data_018_d3;
reg       [7:0] vec_data_019;
reg       [7:0] vec_data_019_d2;
reg       [7:0] vec_data_019_d3;
reg       [7:0] vec_data_020;
reg       [7:0] vec_data_020_d2;
reg       [7:0] vec_data_020_d3;
reg       [7:0] vec_data_021;
reg       [7:0] vec_data_021_d2;
reg       [7:0] vec_data_021_d3;
reg       [7:0] vec_data_022;
reg       [7:0] vec_data_022_d2;
reg       [7:0] vec_data_022_d3;
reg       [7:0] vec_data_023;
reg       [7:0] vec_data_023_d2;
reg       [7:0] vec_data_023_d3;
reg       [7:0] vec_data_024;
reg       [7:0] vec_data_024_d2;
reg       [7:0] vec_data_024_d3;
reg       [7:0] vec_data_025;
reg       [7:0] vec_data_025_d2;
reg       [7:0] vec_data_025_d3;
reg       [7:0] vec_data_026;
reg       [7:0] vec_data_026_d2;
reg       [7:0] vec_data_026_d3;
reg       [7:0] vec_data_027;
reg       [7:0] vec_data_027_d2;
reg       [7:0] vec_data_027_d3;
reg       [7:0] vec_data_028;
reg       [7:0] vec_data_028_d2;
reg       [7:0] vec_data_028_d3;
reg       [7:0] vec_data_029;
reg       [7:0] vec_data_029_d2;
reg       [7:0] vec_data_029_d3;
reg       [7:0] vec_data_030;
reg       [7:0] vec_data_030_d2;
reg       [7:0] vec_data_030_d3;
reg       [7:0] vec_data_031;
reg       [7:0] vec_data_031_d2;
reg       [7:0] vec_data_031_d3;
reg       [7:0] vec_data_032;
reg       [7:0] vec_data_032_d2;
reg       [7:0] vec_data_032_d3;
reg       [7:0] vec_data_033;
reg       [7:0] vec_data_033_d2;
reg       [7:0] vec_data_033_d3;
reg       [7:0] vec_data_034;
reg       [7:0] vec_data_034_d2;
reg       [7:0] vec_data_034_d3;
reg       [7:0] vec_data_035;
reg       [7:0] vec_data_035_d2;
reg       [7:0] vec_data_035_d3;
reg       [7:0] vec_data_036;
reg       [7:0] vec_data_036_d2;
reg       [7:0] vec_data_036_d3;
reg       [7:0] vec_data_037;
reg       [7:0] vec_data_037_d2;
reg       [7:0] vec_data_037_d3;
reg       [7:0] vec_data_038;
reg       [7:0] vec_data_038_d2;
reg       [7:0] vec_data_038_d3;
reg       [7:0] vec_data_039;
reg       [7:0] vec_data_039_d2;
reg       [7:0] vec_data_039_d3;
reg       [7:0] vec_data_040;
reg       [7:0] vec_data_040_d2;
reg       [7:0] vec_data_040_d3;
reg       [7:0] vec_data_041;
reg       [7:0] vec_data_041_d2;
reg       [7:0] vec_data_041_d3;
reg       [7:0] vec_data_042;
reg       [7:0] vec_data_042_d2;
reg       [7:0] vec_data_042_d3;
reg       [7:0] vec_data_043;
reg       [7:0] vec_data_043_d2;
reg       [7:0] vec_data_043_d3;
reg       [7:0] vec_data_044;
reg       [7:0] vec_data_044_d2;
reg       [7:0] vec_data_044_d3;
reg       [7:0] vec_data_045;
reg       [7:0] vec_data_045_d2;
reg       [7:0] vec_data_045_d3;
reg       [7:0] vec_data_046;
reg       [7:0] vec_data_046_d2;
reg       [7:0] vec_data_046_d3;
reg       [7:0] vec_data_047;
reg       [7:0] vec_data_047_d2;
reg       [7:0] vec_data_047_d3;
reg       [7:0] vec_data_048;
reg       [7:0] vec_data_048_d2;
reg       [7:0] vec_data_048_d3;
reg       [7:0] vec_data_049;
reg       [7:0] vec_data_049_d2;
reg       [7:0] vec_data_049_d3;
reg       [7:0] vec_data_050;
reg       [7:0] vec_data_050_d2;
reg       [7:0] vec_data_050_d3;
reg       [7:0] vec_data_051;
reg       [7:0] vec_data_051_d2;
reg       [7:0] vec_data_051_d3;
reg       [7:0] vec_data_052;
reg       [7:0] vec_data_052_d2;
reg       [7:0] vec_data_052_d3;
reg       [7:0] vec_data_053;
reg       [7:0] vec_data_053_d2;
reg       [7:0] vec_data_053_d3;
reg       [7:0] vec_data_054;
reg       [7:0] vec_data_054_d2;
reg       [7:0] vec_data_054_d3;
reg       [7:0] vec_data_055;
reg       [7:0] vec_data_055_d2;
reg       [7:0] vec_data_055_d3;
reg       [7:0] vec_data_056;
reg       [7:0] vec_data_056_d2;
reg       [7:0] vec_data_056_d3;
reg       [7:0] vec_data_057;
reg       [7:0] vec_data_057_d2;
reg       [7:0] vec_data_057_d3;
reg       [7:0] vec_data_058;
reg       [7:0] vec_data_058_d2;
reg       [7:0] vec_data_058_d3;
reg       [7:0] vec_data_059;
reg       [7:0] vec_data_059_d2;
reg       [7:0] vec_data_059_d3;
reg       [7:0] vec_data_060;
reg       [7:0] vec_data_060_d2;
reg       [7:0] vec_data_060_d3;
reg       [7:0] vec_data_061;
reg       [7:0] vec_data_061_d2;
reg       [7:0] vec_data_061_d3;
reg       [7:0] vec_data_062;
reg       [7:0] vec_data_062_d2;
reg       [7:0] vec_data_062_d3;
reg       [7:0] vec_data_063;
reg       [7:0] vec_data_063_d2;
reg       [7:0] vec_data_063_d3;
reg       [7:0] vec_data_064;
reg       [7:0] vec_data_064_d2;
reg       [7:0] vec_data_064_d3;
reg       [7:0] vec_data_065;
reg       [7:0] vec_data_065_d2;
reg       [7:0] vec_data_065_d3;
reg       [7:0] vec_data_066;
reg       [7:0] vec_data_066_d2;
reg       [7:0] vec_data_066_d3;
reg       [7:0] vec_data_067;
reg       [7:0] vec_data_067_d2;
reg       [7:0] vec_data_067_d3;
reg       [7:0] vec_data_068;
reg       [7:0] vec_data_068_d2;
reg       [7:0] vec_data_068_d3;
reg       [7:0] vec_data_069;
reg       [7:0] vec_data_069_d2;
reg       [7:0] vec_data_069_d3;
reg       [7:0] vec_data_070;
reg       [7:0] vec_data_070_d2;
reg       [7:0] vec_data_070_d3;
reg       [7:0] vec_data_071;
reg       [7:0] vec_data_071_d2;
reg       [7:0] vec_data_071_d3;
reg       [7:0] vec_data_072;
reg       [7:0] vec_data_072_d2;
reg       [7:0] vec_data_072_d3;
reg       [7:0] vec_data_073;
reg       [7:0] vec_data_073_d2;
reg       [7:0] vec_data_073_d3;
reg       [7:0] vec_data_074;
reg       [7:0] vec_data_074_d2;
reg       [7:0] vec_data_074_d3;
reg       [7:0] vec_data_075;
reg       [7:0] vec_data_075_d2;
reg       [7:0] vec_data_075_d3;
reg       [7:0] vec_data_076;
reg       [7:0] vec_data_076_d2;
reg       [7:0] vec_data_076_d3;
reg       [7:0] vec_data_077;
reg       [7:0] vec_data_077_d2;
reg       [7:0] vec_data_077_d3;
reg       [7:0] vec_data_078;
reg       [7:0] vec_data_078_d2;
reg       [7:0] vec_data_078_d3;
reg       [7:0] vec_data_079;
reg       [7:0] vec_data_079_d2;
reg       [7:0] vec_data_079_d3;
reg       [7:0] vec_data_080;
reg       [7:0] vec_data_080_d2;
reg       [7:0] vec_data_080_d3;
reg       [7:0] vec_data_081;
reg       [7:0] vec_data_081_d2;
reg       [7:0] vec_data_081_d3;
reg       [7:0] vec_data_082;
reg       [7:0] vec_data_082_d2;
reg       [7:0] vec_data_082_d3;
reg       [7:0] vec_data_083;
reg       [7:0] vec_data_083_d2;
reg       [7:0] vec_data_083_d3;
reg       [7:0] vec_data_084;
reg       [7:0] vec_data_084_d2;
reg       [7:0] vec_data_084_d3;
reg       [7:0] vec_data_085;
reg       [7:0] vec_data_085_d2;
reg       [7:0] vec_data_085_d3;
reg       [7:0] vec_data_086;
reg       [7:0] vec_data_086_d2;
reg       [7:0] vec_data_086_d3;
reg       [7:0] vec_data_087;
reg       [7:0] vec_data_087_d2;
reg       [7:0] vec_data_087_d3;
reg       [7:0] vec_data_088;
reg       [7:0] vec_data_088_d2;
reg       [7:0] vec_data_088_d3;
reg       [7:0] vec_data_089;
reg       [7:0] vec_data_089_d2;
reg       [7:0] vec_data_089_d3;
reg       [7:0] vec_data_090;
reg       [7:0] vec_data_090_d2;
reg       [7:0] vec_data_090_d3;
reg       [7:0] vec_data_091;
reg       [7:0] vec_data_091_d2;
reg       [7:0] vec_data_091_d3;
reg       [7:0] vec_data_092;
reg       [7:0] vec_data_092_d2;
reg       [7:0] vec_data_092_d3;
reg       [7:0] vec_data_093;
reg       [7:0] vec_data_093_d2;
reg       [7:0] vec_data_093_d3;
reg       [7:0] vec_data_094;
reg       [7:0] vec_data_094_d2;
reg       [7:0] vec_data_094_d3;
reg       [7:0] vec_data_095;
reg       [7:0] vec_data_095_d2;
reg       [7:0] vec_data_095_d3;
reg       [7:0] vec_data_096;
reg       [7:0] vec_data_096_d2;
reg       [7:0] vec_data_096_d3;
reg       [7:0] vec_data_097;
reg       [7:0] vec_data_097_d2;
reg       [7:0] vec_data_097_d3;
reg       [7:0] vec_data_098;
reg       [7:0] vec_data_098_d2;
reg       [7:0] vec_data_098_d3;
reg       [7:0] vec_data_099;
reg       [7:0] vec_data_099_d2;
reg       [7:0] vec_data_099_d3;
reg       [7:0] vec_data_100;
reg       [7:0] vec_data_100_d2;
reg       [7:0] vec_data_100_d3;
reg       [7:0] vec_data_101;
reg       [7:0] vec_data_101_d2;
reg       [7:0] vec_data_101_d3;
reg       [7:0] vec_data_102;
reg       [7:0] vec_data_102_d2;
reg       [7:0] vec_data_102_d3;
reg       [7:0] vec_data_103;
reg       [7:0] vec_data_103_d2;
reg       [7:0] vec_data_103_d3;
reg       [7:0] vec_data_104;
reg       [7:0] vec_data_104_d2;
reg       [7:0] vec_data_104_d3;
reg       [7:0] vec_data_105;
reg       [7:0] vec_data_105_d2;
reg       [7:0] vec_data_105_d3;
reg       [7:0] vec_data_106;
reg       [7:0] vec_data_106_d2;
reg       [7:0] vec_data_106_d3;
reg       [7:0] vec_data_107;
reg       [7:0] vec_data_107_d2;
reg       [7:0] vec_data_107_d3;
reg       [7:0] vec_data_108;
reg       [7:0] vec_data_108_d2;
reg       [7:0] vec_data_108_d3;
reg       [7:0] vec_data_109;
reg       [7:0] vec_data_109_d2;
reg       [7:0] vec_data_109_d3;
reg       [7:0] vec_data_110;
reg       [7:0] vec_data_110_d2;
reg       [7:0] vec_data_110_d3;
reg       [7:0] vec_data_111;
reg       [7:0] vec_data_111_d2;
reg       [7:0] vec_data_111_d3;
reg       [7:0] vec_data_112;
reg       [7:0] vec_data_112_d2;
reg       [7:0] vec_data_112_d3;
reg       [7:0] vec_data_113;
reg       [7:0] vec_data_113_d2;
reg       [7:0] vec_data_113_d3;
reg       [7:0] vec_data_114;
reg       [7:0] vec_data_114_d2;
reg       [7:0] vec_data_114_d3;
reg       [7:0] vec_data_115;
reg       [7:0] vec_data_115_d2;
reg       [7:0] vec_data_115_d3;
reg       [7:0] vec_data_116;
reg       [7:0] vec_data_116_d2;
reg       [7:0] vec_data_116_d3;
reg       [7:0] vec_data_117;
reg       [7:0] vec_data_117_d2;
reg       [7:0] vec_data_117_d3;
reg       [7:0] vec_data_118;
reg       [7:0] vec_data_118_d2;
reg       [7:0] vec_data_118_d3;
reg       [7:0] vec_data_119;
reg       [7:0] vec_data_119_d2;
reg       [7:0] vec_data_119_d3;
reg       [7:0] vec_data_120;
reg       [7:0] vec_data_120_d2;
reg       [7:0] vec_data_120_d3;
reg       [7:0] vec_data_121;
reg       [7:0] vec_data_121_d2;
reg       [7:0] vec_data_121_d3;
reg       [7:0] vec_data_122;
reg       [7:0] vec_data_122_d2;
reg       [7:0] vec_data_122_d3;
reg       [7:0] vec_data_123;
reg       [7:0] vec_data_123_d2;
reg       [7:0] vec_data_123_d3;
reg       [7:0] vec_data_124;
reg       [7:0] vec_data_124_d2;
reg       [7:0] vec_data_124_d3;
reg       [7:0] vec_data_125;
reg       [7:0] vec_data_125_d2;
reg       [7:0] vec_data_125_d3;
reg       [7:0] vec_data_126;
reg       [7:0] vec_data_126_d2;
reg       [7:0] vec_data_126_d3;
reg       [7:0] vec_data_127;
reg       [7:0] vec_data_127_d2;
reg       [7:0] vec_data_127_d3;
reg       [0:0] vec_sum_000;
reg             vec_sum_000_d1;
reg       [1:0] vec_sum_001;
reg       [1:0] vec_sum_001_d1;
reg       [1:0] vec_sum_002;
reg       [1:0] vec_sum_002_d1;
reg       [2:0] vec_sum_003;
reg       [2:0] vec_sum_003_d1;
reg       [2:0] vec_sum_004;
reg       [2:0] vec_sum_004_d1;
reg       [2:0] vec_sum_005;
reg       [2:0] vec_sum_005_d1;
reg       [2:0] vec_sum_006;
reg       [2:0] vec_sum_006_d1;
reg       [3:0] vec_sum_007;
reg       [3:0] vec_sum_007_d1;
reg       [3:0] vec_sum_008;
reg       [3:0] vec_sum_008_d1;
reg       [3:0] vec_sum_009;
reg       [3:0] vec_sum_009_d1;
reg       [3:0] vec_sum_010;
reg       [3:0] vec_sum_010_d1;
reg       [3:0] vec_sum_011;
reg       [3:0] vec_sum_011_d1;
reg       [3:0] vec_sum_012;
reg       [3:0] vec_sum_012_d1;
reg       [3:0] vec_sum_013;
reg       [3:0] vec_sum_013_d1;
reg       [3:0] vec_sum_014;
reg       [3:0] vec_sum_014_d1;
reg       [4:0] vec_sum_015;
reg       [4:0] vec_sum_015_d1;
reg       [4:0] vec_sum_016;
reg       [4:0] vec_sum_016_d1;
reg       [4:0] vec_sum_017;
reg       [4:0] vec_sum_017_d1;
reg       [4:0] vec_sum_018;
reg       [4:0] vec_sum_018_d1;
reg       [4:0] vec_sum_019;
reg       [4:0] vec_sum_019_d1;
reg       [4:0] vec_sum_020;
reg       [4:0] vec_sum_020_d1;
reg       [4:0] vec_sum_021;
reg       [4:0] vec_sum_021_d1;
reg       [4:0] vec_sum_022;
reg       [4:0] vec_sum_022_d1;
reg       [4:0] vec_sum_023;
reg       [4:0] vec_sum_023_d1;
reg       [4:0] vec_sum_024;
reg       [4:0] vec_sum_024_d1;
reg       [4:0] vec_sum_025;
reg       [4:0] vec_sum_025_d1;
reg       [4:0] vec_sum_026;
reg       [4:0] vec_sum_026_d1;
reg       [4:0] vec_sum_027;
reg       [4:0] vec_sum_027_d1;
reg       [4:0] vec_sum_028;
reg       [4:0] vec_sum_028_d1;
reg       [4:0] vec_sum_029;
reg       [4:0] vec_sum_029_d1;
reg       [4:0] vec_sum_030;
reg       [4:0] vec_sum_030_d1;
reg       [5:0] vec_sum_031;
reg       [5:0] vec_sum_031_d1;
reg       [5:0] vec_sum_032;
reg       [5:0] vec_sum_032_d1;
reg       [5:0] vec_sum_033;
reg       [5:0] vec_sum_033_d1;
reg       [5:0] vec_sum_034;
reg       [5:0] vec_sum_034_d1;
reg       [5:0] vec_sum_035;
reg       [5:0] vec_sum_035_d1;
reg       [5:0] vec_sum_036;
reg       [5:0] vec_sum_036_d1;
reg       [5:0] vec_sum_037;
reg       [5:0] vec_sum_037_d1;
reg       [5:0] vec_sum_038;
reg       [5:0] vec_sum_038_d1;
reg       [5:0] vec_sum_039;
reg       [5:0] vec_sum_039_d1;
reg       [5:0] vec_sum_040;
reg       [5:0] vec_sum_040_d1;
reg       [5:0] vec_sum_041;
reg       [5:0] vec_sum_041_d1;
reg       [5:0] vec_sum_042;
reg       [5:0] vec_sum_042_d1;
reg       [5:0] vec_sum_043;
reg       [5:0] vec_sum_043_d1;
reg       [5:0] vec_sum_044;
reg       [5:0] vec_sum_044_d1;
reg       [5:0] vec_sum_045;
reg       [5:0] vec_sum_045_d1;
reg       [5:0] vec_sum_046;
reg       [5:0] vec_sum_046_d1;
reg       [5:0] vec_sum_047;
reg       [5:0] vec_sum_047_d1;
reg       [5:0] vec_sum_048;
reg       [5:0] vec_sum_048_d1;
reg       [5:0] vec_sum_049;
reg       [5:0] vec_sum_049_d1;
reg       [5:0] vec_sum_050;
reg       [5:0] vec_sum_050_d1;
reg       [5:0] vec_sum_051;
reg       [5:0] vec_sum_051_d1;
reg       [5:0] vec_sum_052;
reg       [5:0] vec_sum_052_d1;
reg       [5:0] vec_sum_053;
reg       [5:0] vec_sum_053_d1;
reg       [5:0] vec_sum_054;
reg       [5:0] vec_sum_054_d1;
reg       [5:0] vec_sum_055;
reg       [5:0] vec_sum_055_d1;
reg       [5:0] vec_sum_056;
reg       [5:0] vec_sum_056_d1;
reg       [5:0] vec_sum_057;
reg       [5:0] vec_sum_057_d1;
reg       [5:0] vec_sum_058;
reg       [5:0] vec_sum_058_d1;
reg       [5:0] vec_sum_059;
reg       [5:0] vec_sum_059_d1;
reg       [5:0] vec_sum_060;
reg       [5:0] vec_sum_060_d1;
reg       [5:0] vec_sum_061;
reg       [5:0] vec_sum_061_d1;
reg       [5:0] vec_sum_062;
reg       [5:0] vec_sum_062_d1;
reg       [6:0] vec_sum_063;
reg       [6:0] vec_sum_063_d1;
reg       [6:0] vec_sum_064;
reg       [6:0] vec_sum_064_d1;
reg       [6:0] vec_sum_065;
reg       [6:0] vec_sum_065_d1;
reg       [6:0] vec_sum_066;
reg       [6:0] vec_sum_066_d1;
reg       [6:0] vec_sum_067;
reg       [6:0] vec_sum_067_d1;
reg       [6:0] vec_sum_068;
reg       [6:0] vec_sum_068_d1;
reg       [6:0] vec_sum_069;
reg       [6:0] vec_sum_069_d1;
reg       [6:0] vec_sum_070;
reg       [6:0] vec_sum_070_d1;
reg       [6:0] vec_sum_071;
reg       [6:0] vec_sum_071_d1;
reg       [6:0] vec_sum_072;
reg       [6:0] vec_sum_072_d1;
reg       [6:0] vec_sum_073;
reg       [6:0] vec_sum_073_d1;
reg       [6:0] vec_sum_074;
reg       [6:0] vec_sum_074_d1;
reg       [6:0] vec_sum_075;
reg       [6:0] vec_sum_075_d1;
reg       [6:0] vec_sum_076;
reg       [6:0] vec_sum_076_d1;
reg       [6:0] vec_sum_077;
reg       [6:0] vec_sum_077_d1;
reg       [6:0] vec_sum_078;
reg       [6:0] vec_sum_078_d1;
reg       [6:0] vec_sum_079;
reg       [6:0] vec_sum_079_d1;
reg       [6:0] vec_sum_080;
reg       [6:0] vec_sum_080_d1;
reg       [6:0] vec_sum_081;
reg       [6:0] vec_sum_081_d1;
reg       [6:0] vec_sum_082;
reg       [6:0] vec_sum_082_d1;
reg       [6:0] vec_sum_083;
reg       [6:0] vec_sum_083_d1;
reg       [6:0] vec_sum_084;
reg       [6:0] vec_sum_084_d1;
reg       [6:0] vec_sum_085;
reg       [6:0] vec_sum_085_d1;
reg       [6:0] vec_sum_086;
reg       [6:0] vec_sum_086_d1;
reg       [6:0] vec_sum_087;
reg       [6:0] vec_sum_087_d1;
reg       [6:0] vec_sum_088;
reg       [6:0] vec_sum_088_d1;
reg       [6:0] vec_sum_089;
reg       [6:0] vec_sum_089_d1;
reg       [6:0] vec_sum_090;
reg       [6:0] vec_sum_090_d1;
reg       [6:0] vec_sum_091;
reg       [6:0] vec_sum_091_d1;
reg       [6:0] vec_sum_092;
reg       [6:0] vec_sum_092_d1;
reg       [6:0] vec_sum_093;
reg       [6:0] vec_sum_093_d1;
reg       [6:0] vec_sum_094;
reg       [6:0] vec_sum_094_d1;
reg       [6:0] vec_sum_095;
reg       [6:0] vec_sum_095_d1;
reg       [6:0] vec_sum_096;
reg       [6:0] vec_sum_096_d1;
reg       [6:0] vec_sum_097;
reg       [6:0] vec_sum_097_d1;
reg       [6:0] vec_sum_098;
reg       [6:0] vec_sum_098_d1;
reg       [6:0] vec_sum_099;
reg       [6:0] vec_sum_099_d1;
reg       [6:0] vec_sum_100;
reg       [6:0] vec_sum_100_d1;
reg       [6:0] vec_sum_101;
reg       [6:0] vec_sum_101_d1;
reg       [6:0] vec_sum_102;
reg       [6:0] vec_sum_102_d1;
reg       [6:0] vec_sum_103;
reg       [6:0] vec_sum_103_d1;
reg       [6:0] vec_sum_104;
reg       [6:0] vec_sum_104_d1;
reg       [6:0] vec_sum_105;
reg       [6:0] vec_sum_105_d1;
reg       [6:0] vec_sum_106;
reg       [6:0] vec_sum_106_d1;
reg       [6:0] vec_sum_107;
reg       [6:0] vec_sum_107_d1;
reg       [6:0] vec_sum_108;
reg       [6:0] vec_sum_108_d1;
reg       [6:0] vec_sum_109;
reg       [6:0] vec_sum_109_d1;
reg       [6:0] vec_sum_110;
reg       [6:0] vec_sum_110_d1;
reg       [6:0] vec_sum_111;
reg       [6:0] vec_sum_111_d1;
reg       [6:0] vec_sum_112;
reg       [6:0] vec_sum_112_d1;
reg       [6:0] vec_sum_113;
reg       [6:0] vec_sum_113_d1;
reg       [6:0] vec_sum_114;
reg       [6:0] vec_sum_114_d1;
reg       [6:0] vec_sum_115;
reg       [6:0] vec_sum_115_d1;
reg       [6:0] vec_sum_116;
reg       [6:0] vec_sum_116_d1;
reg       [6:0] vec_sum_117;
reg       [6:0] vec_sum_117_d1;
reg       [6:0] vec_sum_118;
reg       [6:0] vec_sum_118_d1;
reg       [6:0] vec_sum_119;
reg       [6:0] vec_sum_119_d1;
reg       [6:0] vec_sum_120;
reg       [6:0] vec_sum_120_d1;
reg       [6:0] vec_sum_121;
reg       [6:0] vec_sum_121_d1;
reg       [6:0] vec_sum_122;
reg       [6:0] vec_sum_122_d1;
reg       [6:0] vec_sum_123;
reg       [6:0] vec_sum_123_d1;
reg       [6:0] vec_sum_124;
reg       [6:0] vec_sum_124_d1;
reg       [6:0] vec_sum_125;
reg       [6:0] vec_sum_125_d1;
reg       [6:0] vec_sum_126;
reg       [6:0] vec_sum_126_d1;
reg       [7:0] vec_sum_127;
reg       [7:0] vec_sum_127_d1;

// synoff nets

// monitor nets

// debug nets

// tie high nets

// tie low nets

// no connect nets

// not all bits used nets

// todo nets

    
/////////////////////////////////////////////////////////////////////////////////////////////
// Decoder of compressed weight                                                  
//
//            data_mask             input_data     mac_sel
//                |                     |            |
//            sums_for_sel           register     register
//                |                     |            |
//                ------------------>  mux        register
//                                      |            |
//                                   output_data  output_sel
//
/////////////////////////////////////////////////////////////////////////////////////////////


////////////////////////////////// phase I: calculate sums for mux //////////////////////////////////


assign input_mask_gated = ~input_mask_en[8] ? 128'b0 : input_mask;

always @(
  input_mask_gated
  ) begin
    vec_sum_000 = input_mask_gated[0];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_001 = input_mask_gated[0] + input_mask_gated[1];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_002 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_003 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_004 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_005 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_006 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_007 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_008 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_009 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_010 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_011 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_012 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_013 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_014 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_015 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_016 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_017 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_018 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_019 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_020 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_021 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_022 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_023 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_024 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_025 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_026 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_027 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_028 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_029 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_030 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_031 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_032 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_033 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_034 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_035 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_036 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_037 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_038 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_039 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_040 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_041 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_042 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_043 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_044 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_045 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_046 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_047 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_048 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_049 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_050 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_051 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_052 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_053 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_054 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_055 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_056 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_057 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_058 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_059 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_060 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_061 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_062 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_063 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_064 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_065 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_066 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_067 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_068 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_069 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_070 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_071 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_072 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_073 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_074 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_075 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_076 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_077 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_078 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_079 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_080 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_081 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_082 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_083 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_084 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_085 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_086 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_087 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_088 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_089 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_090 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_091 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_092 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_093 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_094 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_095 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_096 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_097 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_098 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_099 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_100 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_101 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_102 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_103 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_104 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_105 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_106 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_107 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_108 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_109 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_110 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_111 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_112 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_113 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_114 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_115 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_116 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_117 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_118 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_119 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_120 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_121 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_122 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121] + input_mask_gated[122];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_123 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121] + input_mask_gated[122] + input_mask_gated[123];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_124 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121] + input_mask_gated[122] + input_mask_gated[123] + input_mask_gated[124];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_125 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121] + input_mask_gated[122] + input_mask_gated[123] + input_mask_gated[124] + input_mask_gated[125];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_126 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121] + input_mask_gated[122] + input_mask_gated[123] + input_mask_gated[124] + input_mask_gated[125] + input_mask_gated[126];
end

always @(
  input_mask_gated
  ) begin
    vec_sum_127 = input_mask_gated[0] + input_mask_gated[1] + input_mask_gated[2] + input_mask_gated[3] + input_mask_gated[4] + input_mask_gated[5] + input_mask_gated[6] + input_mask_gated[7]
                + input_mask_gated[8] + input_mask_gated[9] + input_mask_gated[10] + input_mask_gated[11] + input_mask_gated[12] + input_mask_gated[13] + input_mask_gated[14] + input_mask_gated[15]
                + input_mask_gated[16] + input_mask_gated[17] + input_mask_gated[18] + input_mask_gated[19] + input_mask_gated[20] + input_mask_gated[21] + input_mask_gated[22] + input_mask_gated[23]
                + input_mask_gated[24] + input_mask_gated[25] + input_mask_gated[26] + input_mask_gated[27] + input_mask_gated[28] + input_mask_gated[29] + input_mask_gated[30] + input_mask_gated[31]
                + input_mask_gated[32] + input_mask_gated[33] + input_mask_gated[34] + input_mask_gated[35] + input_mask_gated[36] + input_mask_gated[37] + input_mask_gated[38] + input_mask_gated[39]
                + input_mask_gated[40] + input_mask_gated[41] + input_mask_gated[42] + input_mask_gated[43] + input_mask_gated[44] + input_mask_gated[45] + input_mask_gated[46] + input_mask_gated[47]
                + input_mask_gated[48] + input_mask_gated[49] + input_mask_gated[50] + input_mask_gated[51] + input_mask_gated[52] + input_mask_gated[53] + input_mask_gated[54] + input_mask_gated[55]
                + input_mask_gated[56] + input_mask_gated[57] + input_mask_gated[58] + input_mask_gated[59] + input_mask_gated[60] + input_mask_gated[61] + input_mask_gated[62] + input_mask_gated[63]
                + input_mask_gated[64] + input_mask_gated[65] + input_mask_gated[66] + input_mask_gated[67] + input_mask_gated[68] + input_mask_gated[69] + input_mask_gated[70] + input_mask_gated[71]
                + input_mask_gated[72] + input_mask_gated[73] + input_mask_gated[74] + input_mask_gated[75] + input_mask_gated[76] + input_mask_gated[77] + input_mask_gated[78] + input_mask_gated[79]
                + input_mask_gated[80] + input_mask_gated[81] + input_mask_gated[82] + input_mask_gated[83] + input_mask_gated[84] + input_mask_gated[85] + input_mask_gated[86] + input_mask_gated[87]
                + input_mask_gated[88] + input_mask_gated[89] + input_mask_gated[90] + input_mask_gated[91] + input_mask_gated[92] + input_mask_gated[93] + input_mask_gated[94] + input_mask_gated[95]
                + input_mask_gated[96] + input_mask_gated[97] + input_mask_gated[98] + input_mask_gated[99] + input_mask_gated[100] + input_mask_gated[101] + input_mask_gated[102] + input_mask_gated[103]
                + input_mask_gated[104] + input_mask_gated[105] + input_mask_gated[106] + input_mask_gated[107] + input_mask_gated[108] + input_mask_gated[109] + input_mask_gated[110] + input_mask_gated[111]
                + input_mask_gated[112] + input_mask_gated[113] + input_mask_gated[114] + input_mask_gated[115] + input_mask_gated[116] + input_mask_gated[117] + input_mask_gated[118] + input_mask_gated[119]
                + input_mask_gated[120] + input_mask_gated[121] + input_mask_gated[122] + input_mask_gated[123] + input_mask_gated[124] + input_mask_gated[125] + input_mask_gated[126] + input_mask_gated[127];
end



////////////////////////////////// phase I: registers //////////////////////////////////
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    valid_d1 <= 1'b0;
  end else begin
  valid_d1 <= input_pipe_valid;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid) == 1'b1) begin
    data_d1 <= input_data;
  // VCS coverage off
  end else if ((input_pipe_valid) == 1'b0) begin
  end else begin
    data_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_mask_en[9]) == 1'b1) begin
    mask_d1 <= input_mask;
  // VCS coverage off
  end else if ((input_mask_en[9]) == 1'b0) begin
  end else begin
    mask_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid) == 1'b1) begin
    sel_d1 <= input_sel;
  // VCS coverage off
  end else if ((input_pipe_valid) == 1'b0) begin
  end else begin
    sel_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_000_d1 <= vec_sum_000;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_000_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_001_d1 <= vec_sum_001;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_001_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_002_d1 <= vec_sum_002;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_002_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_003_d1 <= vec_sum_003;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_003_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_004_d1 <= vec_sum_004;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_004_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_005_d1 <= vec_sum_005;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_005_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_006_d1 <= vec_sum_006;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_006_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_007_d1 <= vec_sum_007;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_007_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_008_d1 <= vec_sum_008;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_008_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_009_d1 <= vec_sum_009;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_009_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_010_d1 <= vec_sum_010;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_010_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_011_d1 <= vec_sum_011;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_011_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_012_d1 <= vec_sum_012;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_012_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_013_d1 <= vec_sum_013;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_013_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_014_d1 <= vec_sum_014;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_014_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[0]) == 1'b1) begin
    vec_sum_015_d1 <= vec_sum_015;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[0]) == 1'b0) begin
  end else begin
    vec_sum_015_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_016_d1 <= vec_sum_016;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_016_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_017_d1 <= vec_sum_017;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_017_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_018_d1 <= vec_sum_018;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_018_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_019_d1 <= vec_sum_019;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_019_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_020_d1 <= vec_sum_020;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_020_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_021_d1 <= vec_sum_021;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_021_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_022_d1 <= vec_sum_022;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_022_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_023_d1 <= vec_sum_023;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_023_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_024_d1 <= vec_sum_024;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_024_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_025_d1 <= vec_sum_025;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_025_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_026_d1 <= vec_sum_026;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_026_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_027_d1 <= vec_sum_027;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_027_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_028_d1 <= vec_sum_028;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_028_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_029_d1 <= vec_sum_029;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_029_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_030_d1 <= vec_sum_030;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_030_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[1]) == 1'b1) begin
    vec_sum_031_d1 <= vec_sum_031;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[1]) == 1'b0) begin
  end else begin
    vec_sum_031_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_032_d1 <= vec_sum_032;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_032_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_033_d1 <= vec_sum_033;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_033_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_034_d1 <= vec_sum_034;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_034_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_035_d1 <= vec_sum_035;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_035_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_036_d1 <= vec_sum_036;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_036_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_037_d1 <= vec_sum_037;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_037_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_038_d1 <= vec_sum_038;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_038_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_039_d1 <= vec_sum_039;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_039_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_040_d1 <= vec_sum_040;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_040_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_041_d1 <= vec_sum_041;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_041_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_042_d1 <= vec_sum_042;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_042_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_043_d1 <= vec_sum_043;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_043_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_044_d1 <= vec_sum_044;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_044_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_045_d1 <= vec_sum_045;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_045_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_046_d1 <= vec_sum_046;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_046_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[2]) == 1'b1) begin
    vec_sum_047_d1 <= vec_sum_047;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[2]) == 1'b0) begin
  end else begin
    vec_sum_047_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_048_d1 <= vec_sum_048;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_048_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_049_d1 <= vec_sum_049;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_049_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_050_d1 <= vec_sum_050;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_050_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_051_d1 <= vec_sum_051;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_051_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_052_d1 <= vec_sum_052;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_052_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_053_d1 <= vec_sum_053;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_053_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_054_d1 <= vec_sum_054;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_054_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_055_d1 <= vec_sum_055;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_055_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_056_d1 <= vec_sum_056;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_056_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_057_d1 <= vec_sum_057;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_057_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_058_d1 <= vec_sum_058;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_058_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_059_d1 <= vec_sum_059;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_059_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_060_d1 <= vec_sum_060;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_060_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_061_d1 <= vec_sum_061;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_061_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_062_d1 <= vec_sum_062;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_062_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[3]) == 1'b1) begin
    vec_sum_063_d1 <= vec_sum_063;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[3]) == 1'b0) begin
  end else begin
    vec_sum_063_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_064_d1 <= vec_sum_064;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_064_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_065_d1 <= vec_sum_065;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_065_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_066_d1 <= vec_sum_066;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_066_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_067_d1 <= vec_sum_067;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_067_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_068_d1 <= vec_sum_068;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_068_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_069_d1 <= vec_sum_069;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_069_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_070_d1 <= vec_sum_070;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_070_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_071_d1 <= vec_sum_071;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_071_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_072_d1 <= vec_sum_072;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_072_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_073_d1 <= vec_sum_073;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_073_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_074_d1 <= vec_sum_074;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_074_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_075_d1 <= vec_sum_075;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_075_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_076_d1 <= vec_sum_076;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_076_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_077_d1 <= vec_sum_077;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_077_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_078_d1 <= vec_sum_078;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_078_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[4]) == 1'b1) begin
    vec_sum_079_d1 <= vec_sum_079;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[4]) == 1'b0) begin
  end else begin
    vec_sum_079_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_080_d1 <= vec_sum_080;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_080_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_081_d1 <= vec_sum_081;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_081_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_082_d1 <= vec_sum_082;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_082_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_083_d1 <= vec_sum_083;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_083_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_084_d1 <= vec_sum_084;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_084_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_085_d1 <= vec_sum_085;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_085_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_086_d1 <= vec_sum_086;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_086_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_087_d1 <= vec_sum_087;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_087_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_088_d1 <= vec_sum_088;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_088_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_089_d1 <= vec_sum_089;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_089_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_090_d1 <= vec_sum_090;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_090_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_091_d1 <= vec_sum_091;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_091_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_092_d1 <= vec_sum_092;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_092_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_093_d1 <= vec_sum_093;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_093_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_094_d1 <= vec_sum_094;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_094_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[5]) == 1'b1) begin
    vec_sum_095_d1 <= vec_sum_095;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[5]) == 1'b0) begin
  end else begin
    vec_sum_095_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_096_d1 <= vec_sum_096;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_096_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_097_d1 <= vec_sum_097;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_097_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_098_d1 <= vec_sum_098;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_098_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_099_d1 <= vec_sum_099;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_099_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_100_d1 <= vec_sum_100;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_100_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_101_d1 <= vec_sum_101;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_101_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_102_d1 <= vec_sum_102;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_102_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_103_d1 <= vec_sum_103;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_103_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_104_d1 <= vec_sum_104;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_104_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_105_d1 <= vec_sum_105;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_105_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_106_d1 <= vec_sum_106;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_106_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_107_d1 <= vec_sum_107;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_107_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_108_d1 <= vec_sum_108;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_108_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_109_d1 <= vec_sum_109;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_109_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_110_d1 <= vec_sum_110;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_110_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[6]) == 1'b1) begin
    vec_sum_111_d1 <= vec_sum_111;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[6]) == 1'b0) begin
  end else begin
    vec_sum_111_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_112_d1 <= vec_sum_112;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_112_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_113_d1 <= vec_sum_113;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_113_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_114_d1 <= vec_sum_114;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_114_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_115_d1 <= vec_sum_115;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_115_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_116_d1 <= vec_sum_116;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_116_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_117_d1 <= vec_sum_117;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_117_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_118_d1 <= vec_sum_118;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_118_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_119_d1 <= vec_sum_119;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_119_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_120_d1 <= vec_sum_120;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_120_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_121_d1 <= vec_sum_121;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_121_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_122_d1 <= vec_sum_122;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_122_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_123_d1 <= vec_sum_123;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_123_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_124_d1 <= vec_sum_124;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_124_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_125_d1 <= vec_sum_125;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_125_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_126_d1 <= vec_sum_126;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_126_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((input_pipe_valid & input_mask_en[7]) == 1'b1) begin
    vec_sum_127_d1 <= vec_sum_127;
  // VCS coverage off
  end else if ((input_pipe_valid & input_mask_en[7]) == 1'b0) begin
  end else begin
    vec_sum_127_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


////////////////////////////////// phase II: mux //////////////////////////////////
always @(
  vec_sum_000_d1
  or data_d1
  ) begin
    vec_data_000 = 8'b0;
    case(vec_sum_000_d1)
        1'd1: vec_data_000 = data_d1[7:0];
    endcase
end

always @(
  vec_sum_001_d1
  or data_d1
  ) begin
    vec_data_001 = 8'b0;
    case(vec_sum_001_d1)
        2'd1: vec_data_001 = data_d1[7:0];
        2'd2: vec_data_001 = data_d1[15:8];
    endcase
end

always @(
  vec_sum_002_d1
  or data_d1
  ) begin
    vec_data_002 = 8'b0;
    case(vec_sum_002_d1)
        2'd1: vec_data_002 = data_d1[7:0];
        2'd2: vec_data_002 = data_d1[15:8];
        2'd3: vec_data_002 = data_d1[23:16];
    endcase
end

always @(
  vec_sum_003_d1
  or data_d1
  ) begin
    vec_data_003 = 8'b0;
    case(vec_sum_003_d1)
        3'd1: vec_data_003 = data_d1[7:0];
        3'd2: vec_data_003 = data_d1[15:8];
        3'd3: vec_data_003 = data_d1[23:16];
        3'd4: vec_data_003 = data_d1[31:24];
    endcase
end

always @(
  vec_sum_004_d1
  or data_d1
  ) begin
    vec_data_004 = 8'b0;
    case(vec_sum_004_d1)
        3'd1: vec_data_004 = data_d1[7:0];
        3'd2: vec_data_004 = data_d1[15:8];
        3'd3: vec_data_004 = data_d1[23:16];
        3'd4: vec_data_004 = data_d1[31:24];
        3'd5: vec_data_004 = data_d1[39:32];
    endcase
end

always @(
  vec_sum_005_d1
  or data_d1
  ) begin
    vec_data_005 = 8'b0;
    case(vec_sum_005_d1)
        3'd1: vec_data_005 = data_d1[7:0];
        3'd2: vec_data_005 = data_d1[15:8];
        3'd3: vec_data_005 = data_d1[23:16];
        3'd4: vec_data_005 = data_d1[31:24];
        3'd5: vec_data_005 = data_d1[39:32];
        3'd6: vec_data_005 = data_d1[47:40];
    endcase
end

always @(
  vec_sum_006_d1
  or data_d1
  ) begin
    vec_data_006 = 8'b0;
    case(vec_sum_006_d1)
        3'd1: vec_data_006 = data_d1[7:0];
        3'd2: vec_data_006 = data_d1[15:8];
        3'd3: vec_data_006 = data_d1[23:16];
        3'd4: vec_data_006 = data_d1[31:24];
        3'd5: vec_data_006 = data_d1[39:32];
        3'd6: vec_data_006 = data_d1[47:40];
        3'd7: vec_data_006 = data_d1[55:48];
    endcase
end

always @(
  vec_sum_007_d1
  or data_d1
  ) begin
    vec_data_007 = 8'b0;
    case(vec_sum_007_d1)
        4'd1: vec_data_007 = data_d1[7:0];
        4'd2: vec_data_007 = data_d1[15:8];
        4'd3: vec_data_007 = data_d1[23:16];
        4'd4: vec_data_007 = data_d1[31:24];
        4'd5: vec_data_007 = data_d1[39:32];
        4'd6: vec_data_007 = data_d1[47:40];
        4'd7: vec_data_007 = data_d1[55:48];
        4'd8: vec_data_007 = data_d1[63:56];
    endcase
end

always @(
  vec_sum_008_d1
  or data_d1
  ) begin
    vec_data_008 = 8'b0;
    case(vec_sum_008_d1)
        4'd1: vec_data_008 = data_d1[7:0];
        4'd2: vec_data_008 = data_d1[15:8];
        4'd3: vec_data_008 = data_d1[23:16];
        4'd4: vec_data_008 = data_d1[31:24];
        4'd5: vec_data_008 = data_d1[39:32];
        4'd6: vec_data_008 = data_d1[47:40];
        4'd7: vec_data_008 = data_d1[55:48];
        4'd8: vec_data_008 = data_d1[63:56];
        4'd9: vec_data_008 = data_d1[71:64];
    endcase
end

always @(
  vec_sum_009_d1
  or data_d1
  ) begin
    vec_data_009 = 8'b0;
    case(vec_sum_009_d1)
        4'd1: vec_data_009 = data_d1[7:0];
        4'd2: vec_data_009 = data_d1[15:8];
        4'd3: vec_data_009 = data_d1[23:16];
        4'd4: vec_data_009 = data_d1[31:24];
        4'd5: vec_data_009 = data_d1[39:32];
        4'd6: vec_data_009 = data_d1[47:40];
        4'd7: vec_data_009 = data_d1[55:48];
        4'd8: vec_data_009 = data_d1[63:56];
        4'd9: vec_data_009 = data_d1[71:64];
        4'd10: vec_data_009 = data_d1[79:72];
    endcase
end

always @(
  vec_sum_010_d1
  or data_d1
  ) begin
    vec_data_010 = 8'b0;
    case(vec_sum_010_d1)
        4'd1: vec_data_010 = data_d1[7:0];
        4'd2: vec_data_010 = data_d1[15:8];
        4'd3: vec_data_010 = data_d1[23:16];
        4'd4: vec_data_010 = data_d1[31:24];
        4'd5: vec_data_010 = data_d1[39:32];
        4'd6: vec_data_010 = data_d1[47:40];
        4'd7: vec_data_010 = data_d1[55:48];
        4'd8: vec_data_010 = data_d1[63:56];
        4'd9: vec_data_010 = data_d1[71:64];
        4'd10: vec_data_010 = data_d1[79:72];
        4'd11: vec_data_010 = data_d1[87:80];
    endcase
end

always @(
  vec_sum_011_d1
  or data_d1
  ) begin
    vec_data_011 = 8'b0;
    case(vec_sum_011_d1)
        4'd1: vec_data_011 = data_d1[7:0];
        4'd2: vec_data_011 = data_d1[15:8];
        4'd3: vec_data_011 = data_d1[23:16];
        4'd4: vec_data_011 = data_d1[31:24];
        4'd5: vec_data_011 = data_d1[39:32];
        4'd6: vec_data_011 = data_d1[47:40];
        4'd7: vec_data_011 = data_d1[55:48];
        4'd8: vec_data_011 = data_d1[63:56];
        4'd9: vec_data_011 = data_d1[71:64];
        4'd10: vec_data_011 = data_d1[79:72];
        4'd11: vec_data_011 = data_d1[87:80];
        4'd12: vec_data_011 = data_d1[95:88];
    endcase
end

always @(
  vec_sum_012_d1
  or data_d1
  ) begin
    vec_data_012 = 8'b0;
    case(vec_sum_012_d1)
        4'd1: vec_data_012 = data_d1[7:0];
        4'd2: vec_data_012 = data_d1[15:8];
        4'd3: vec_data_012 = data_d1[23:16];
        4'd4: vec_data_012 = data_d1[31:24];
        4'd5: vec_data_012 = data_d1[39:32];
        4'd6: vec_data_012 = data_d1[47:40];
        4'd7: vec_data_012 = data_d1[55:48];
        4'd8: vec_data_012 = data_d1[63:56];
        4'd9: vec_data_012 = data_d1[71:64];
        4'd10: vec_data_012 = data_d1[79:72];
        4'd11: vec_data_012 = data_d1[87:80];
        4'd12: vec_data_012 = data_d1[95:88];
        4'd13: vec_data_012 = data_d1[103:96];
    endcase
end

always @(
  vec_sum_013_d1
  or data_d1
  ) begin
    vec_data_013 = 8'b0;
    case(vec_sum_013_d1)
        4'd1: vec_data_013 = data_d1[7:0];
        4'd2: vec_data_013 = data_d1[15:8];
        4'd3: vec_data_013 = data_d1[23:16];
        4'd4: vec_data_013 = data_d1[31:24];
        4'd5: vec_data_013 = data_d1[39:32];
        4'd6: vec_data_013 = data_d1[47:40];
        4'd7: vec_data_013 = data_d1[55:48];
        4'd8: vec_data_013 = data_d1[63:56];
        4'd9: vec_data_013 = data_d1[71:64];
        4'd10: vec_data_013 = data_d1[79:72];
        4'd11: vec_data_013 = data_d1[87:80];
        4'd12: vec_data_013 = data_d1[95:88];
        4'd13: vec_data_013 = data_d1[103:96];
        4'd14: vec_data_013 = data_d1[111:104];
    endcase
end

always @(
  vec_sum_014_d1
  or data_d1
  ) begin
    vec_data_014 = 8'b0;
    case(vec_sum_014_d1)
        4'd1: vec_data_014 = data_d1[7:0];
        4'd2: vec_data_014 = data_d1[15:8];
        4'd3: vec_data_014 = data_d1[23:16];
        4'd4: vec_data_014 = data_d1[31:24];
        4'd5: vec_data_014 = data_d1[39:32];
        4'd6: vec_data_014 = data_d1[47:40];
        4'd7: vec_data_014 = data_d1[55:48];
        4'd8: vec_data_014 = data_d1[63:56];
        4'd9: vec_data_014 = data_d1[71:64];
        4'd10: vec_data_014 = data_d1[79:72];
        4'd11: vec_data_014 = data_d1[87:80];
        4'd12: vec_data_014 = data_d1[95:88];
        4'd13: vec_data_014 = data_d1[103:96];
        4'd14: vec_data_014 = data_d1[111:104];
        4'd15: vec_data_014 = data_d1[119:112];
    endcase
end

always @(
  vec_sum_015_d1
  or data_d1
  ) begin
    vec_data_015 = 8'b0;
    case(vec_sum_015_d1)
        5'd1: vec_data_015 = data_d1[7:0];
        5'd2: vec_data_015 = data_d1[15:8];
        5'd3: vec_data_015 = data_d1[23:16];
        5'd4: vec_data_015 = data_d1[31:24];
        5'd5: vec_data_015 = data_d1[39:32];
        5'd6: vec_data_015 = data_d1[47:40];
        5'd7: vec_data_015 = data_d1[55:48];
        5'd8: vec_data_015 = data_d1[63:56];
        5'd9: vec_data_015 = data_d1[71:64];
        5'd10: vec_data_015 = data_d1[79:72];
        5'd11: vec_data_015 = data_d1[87:80];
        5'd12: vec_data_015 = data_d1[95:88];
        5'd13: vec_data_015 = data_d1[103:96];
        5'd14: vec_data_015 = data_d1[111:104];
        5'd15: vec_data_015 = data_d1[119:112];
        5'd16: vec_data_015 = data_d1[127:120];
    endcase
end

always @(
  vec_sum_016_d1
  or data_d1
  ) begin
    vec_data_016 = 8'b0;
    case(vec_sum_016_d1)
        5'd1: vec_data_016 = data_d1[7:0];
        5'd2: vec_data_016 = data_d1[15:8];
        5'd3: vec_data_016 = data_d1[23:16];
        5'd4: vec_data_016 = data_d1[31:24];
        5'd5: vec_data_016 = data_d1[39:32];
        5'd6: vec_data_016 = data_d1[47:40];
        5'd7: vec_data_016 = data_d1[55:48];
        5'd8: vec_data_016 = data_d1[63:56];
        5'd9: vec_data_016 = data_d1[71:64];
        5'd10: vec_data_016 = data_d1[79:72];
        5'd11: vec_data_016 = data_d1[87:80];
        5'd12: vec_data_016 = data_d1[95:88];
        5'd13: vec_data_016 = data_d1[103:96];
        5'd14: vec_data_016 = data_d1[111:104];
        5'd15: vec_data_016 = data_d1[119:112];
        5'd16: vec_data_016 = data_d1[127:120];
        5'd17: vec_data_016 = data_d1[135:128];
    endcase
end

always @(
  vec_sum_017_d1
  or data_d1
  ) begin
    vec_data_017 = 8'b0;
    case(vec_sum_017_d1)
        5'd1: vec_data_017 = data_d1[7:0];
        5'd2: vec_data_017 = data_d1[15:8];
        5'd3: vec_data_017 = data_d1[23:16];
        5'd4: vec_data_017 = data_d1[31:24];
        5'd5: vec_data_017 = data_d1[39:32];
        5'd6: vec_data_017 = data_d1[47:40];
        5'd7: vec_data_017 = data_d1[55:48];
        5'd8: vec_data_017 = data_d1[63:56];
        5'd9: vec_data_017 = data_d1[71:64];
        5'd10: vec_data_017 = data_d1[79:72];
        5'd11: vec_data_017 = data_d1[87:80];
        5'd12: vec_data_017 = data_d1[95:88];
        5'd13: vec_data_017 = data_d1[103:96];
        5'd14: vec_data_017 = data_d1[111:104];
        5'd15: vec_data_017 = data_d1[119:112];
        5'd16: vec_data_017 = data_d1[127:120];
        5'd17: vec_data_017 = data_d1[135:128];
        5'd18: vec_data_017 = data_d1[143:136];
    endcase
end

always @(
  vec_sum_018_d1
  or data_d1
  ) begin
    vec_data_018 = 8'b0;
    case(vec_sum_018_d1)
        5'd1: vec_data_018 = data_d1[7:0];
        5'd2: vec_data_018 = data_d1[15:8];
        5'd3: vec_data_018 = data_d1[23:16];
        5'd4: vec_data_018 = data_d1[31:24];
        5'd5: vec_data_018 = data_d1[39:32];
        5'd6: vec_data_018 = data_d1[47:40];
        5'd7: vec_data_018 = data_d1[55:48];
        5'd8: vec_data_018 = data_d1[63:56];
        5'd9: vec_data_018 = data_d1[71:64];
        5'd10: vec_data_018 = data_d1[79:72];
        5'd11: vec_data_018 = data_d1[87:80];
        5'd12: vec_data_018 = data_d1[95:88];
        5'd13: vec_data_018 = data_d1[103:96];
        5'd14: vec_data_018 = data_d1[111:104];
        5'd15: vec_data_018 = data_d1[119:112];
        5'd16: vec_data_018 = data_d1[127:120];
        5'd17: vec_data_018 = data_d1[135:128];
        5'd18: vec_data_018 = data_d1[143:136];
        5'd19: vec_data_018 = data_d1[151:144];
    endcase
end

always @(
  vec_sum_019_d1
  or data_d1
  ) begin
    vec_data_019 = 8'b0;
    case(vec_sum_019_d1)
        5'd1: vec_data_019 = data_d1[7:0];
        5'd2: vec_data_019 = data_d1[15:8];
        5'd3: vec_data_019 = data_d1[23:16];
        5'd4: vec_data_019 = data_d1[31:24];
        5'd5: vec_data_019 = data_d1[39:32];
        5'd6: vec_data_019 = data_d1[47:40];
        5'd7: vec_data_019 = data_d1[55:48];
        5'd8: vec_data_019 = data_d1[63:56];
        5'd9: vec_data_019 = data_d1[71:64];
        5'd10: vec_data_019 = data_d1[79:72];
        5'd11: vec_data_019 = data_d1[87:80];
        5'd12: vec_data_019 = data_d1[95:88];
        5'd13: vec_data_019 = data_d1[103:96];
        5'd14: vec_data_019 = data_d1[111:104];
        5'd15: vec_data_019 = data_d1[119:112];
        5'd16: vec_data_019 = data_d1[127:120];
        5'd17: vec_data_019 = data_d1[135:128];
        5'd18: vec_data_019 = data_d1[143:136];
        5'd19: vec_data_019 = data_d1[151:144];
        5'd20: vec_data_019 = data_d1[159:152];
    endcase
end

always @(
  vec_sum_020_d1
  or data_d1
  ) begin
    vec_data_020 = 8'b0;
    case(vec_sum_020_d1)
        5'd1: vec_data_020 = data_d1[7:0];
        5'd2: vec_data_020 = data_d1[15:8];
        5'd3: vec_data_020 = data_d1[23:16];
        5'd4: vec_data_020 = data_d1[31:24];
        5'd5: vec_data_020 = data_d1[39:32];
        5'd6: vec_data_020 = data_d1[47:40];
        5'd7: vec_data_020 = data_d1[55:48];
        5'd8: vec_data_020 = data_d1[63:56];
        5'd9: vec_data_020 = data_d1[71:64];
        5'd10: vec_data_020 = data_d1[79:72];
        5'd11: vec_data_020 = data_d1[87:80];
        5'd12: vec_data_020 = data_d1[95:88];
        5'd13: vec_data_020 = data_d1[103:96];
        5'd14: vec_data_020 = data_d1[111:104];
        5'd15: vec_data_020 = data_d1[119:112];
        5'd16: vec_data_020 = data_d1[127:120];
        5'd17: vec_data_020 = data_d1[135:128];
        5'd18: vec_data_020 = data_d1[143:136];
        5'd19: vec_data_020 = data_d1[151:144];
        5'd20: vec_data_020 = data_d1[159:152];
        5'd21: vec_data_020 = data_d1[167:160];
    endcase
end

always @(
  vec_sum_021_d1
  or data_d1
  ) begin
    vec_data_021 = 8'b0;
    case(vec_sum_021_d1)
        5'd1: vec_data_021 = data_d1[7:0];
        5'd2: vec_data_021 = data_d1[15:8];
        5'd3: vec_data_021 = data_d1[23:16];
        5'd4: vec_data_021 = data_d1[31:24];
        5'd5: vec_data_021 = data_d1[39:32];
        5'd6: vec_data_021 = data_d1[47:40];
        5'd7: vec_data_021 = data_d1[55:48];
        5'd8: vec_data_021 = data_d1[63:56];
        5'd9: vec_data_021 = data_d1[71:64];
        5'd10: vec_data_021 = data_d1[79:72];
        5'd11: vec_data_021 = data_d1[87:80];
        5'd12: vec_data_021 = data_d1[95:88];
        5'd13: vec_data_021 = data_d1[103:96];
        5'd14: vec_data_021 = data_d1[111:104];
        5'd15: vec_data_021 = data_d1[119:112];
        5'd16: vec_data_021 = data_d1[127:120];
        5'd17: vec_data_021 = data_d1[135:128];
        5'd18: vec_data_021 = data_d1[143:136];
        5'd19: vec_data_021 = data_d1[151:144];
        5'd20: vec_data_021 = data_d1[159:152];
        5'd21: vec_data_021 = data_d1[167:160];
        5'd22: vec_data_021 = data_d1[175:168];
    endcase
end

always @(
  vec_sum_022_d1
  or data_d1
  ) begin
    vec_data_022 = 8'b0;
    case(vec_sum_022_d1)
        5'd1: vec_data_022 = data_d1[7:0];
        5'd2: vec_data_022 = data_d1[15:8];
        5'd3: vec_data_022 = data_d1[23:16];
        5'd4: vec_data_022 = data_d1[31:24];
        5'd5: vec_data_022 = data_d1[39:32];
        5'd6: vec_data_022 = data_d1[47:40];
        5'd7: vec_data_022 = data_d1[55:48];
        5'd8: vec_data_022 = data_d1[63:56];
        5'd9: vec_data_022 = data_d1[71:64];
        5'd10: vec_data_022 = data_d1[79:72];
        5'd11: vec_data_022 = data_d1[87:80];
        5'd12: vec_data_022 = data_d1[95:88];
        5'd13: vec_data_022 = data_d1[103:96];
        5'd14: vec_data_022 = data_d1[111:104];
        5'd15: vec_data_022 = data_d1[119:112];
        5'd16: vec_data_022 = data_d1[127:120];
        5'd17: vec_data_022 = data_d1[135:128];
        5'd18: vec_data_022 = data_d1[143:136];
        5'd19: vec_data_022 = data_d1[151:144];
        5'd20: vec_data_022 = data_d1[159:152];
        5'd21: vec_data_022 = data_d1[167:160];
        5'd22: vec_data_022 = data_d1[175:168];
        5'd23: vec_data_022 = data_d1[183:176];
    endcase
end

always @(
  vec_sum_023_d1
  or data_d1
  ) begin
    vec_data_023 = 8'b0;
    case(vec_sum_023_d1)
        5'd1: vec_data_023 = data_d1[7:0];
        5'd2: vec_data_023 = data_d1[15:8];
        5'd3: vec_data_023 = data_d1[23:16];
        5'd4: vec_data_023 = data_d1[31:24];
        5'd5: vec_data_023 = data_d1[39:32];
        5'd6: vec_data_023 = data_d1[47:40];
        5'd7: vec_data_023 = data_d1[55:48];
        5'd8: vec_data_023 = data_d1[63:56];
        5'd9: vec_data_023 = data_d1[71:64];
        5'd10: vec_data_023 = data_d1[79:72];
        5'd11: vec_data_023 = data_d1[87:80];
        5'd12: vec_data_023 = data_d1[95:88];
        5'd13: vec_data_023 = data_d1[103:96];
        5'd14: vec_data_023 = data_d1[111:104];
        5'd15: vec_data_023 = data_d1[119:112];
        5'd16: vec_data_023 = data_d1[127:120];
        5'd17: vec_data_023 = data_d1[135:128];
        5'd18: vec_data_023 = data_d1[143:136];
        5'd19: vec_data_023 = data_d1[151:144];
        5'd20: vec_data_023 = data_d1[159:152];
        5'd21: vec_data_023 = data_d1[167:160];
        5'd22: vec_data_023 = data_d1[175:168];
        5'd23: vec_data_023 = data_d1[183:176];
        5'd24: vec_data_023 = data_d1[191:184];
    endcase
end

always @(
  vec_sum_024_d1
  or data_d1
  ) begin
    vec_data_024 = 8'b0;
    case(vec_sum_024_d1)
        5'd1: vec_data_024 = data_d1[7:0];
        5'd2: vec_data_024 = data_d1[15:8];
        5'd3: vec_data_024 = data_d1[23:16];
        5'd4: vec_data_024 = data_d1[31:24];
        5'd5: vec_data_024 = data_d1[39:32];
        5'd6: vec_data_024 = data_d1[47:40];
        5'd7: vec_data_024 = data_d1[55:48];
        5'd8: vec_data_024 = data_d1[63:56];
        5'd9: vec_data_024 = data_d1[71:64];
        5'd10: vec_data_024 = data_d1[79:72];
        5'd11: vec_data_024 = data_d1[87:80];
        5'd12: vec_data_024 = data_d1[95:88];
        5'd13: vec_data_024 = data_d1[103:96];
        5'd14: vec_data_024 = data_d1[111:104];
        5'd15: vec_data_024 = data_d1[119:112];
        5'd16: vec_data_024 = data_d1[127:120];
        5'd17: vec_data_024 = data_d1[135:128];
        5'd18: vec_data_024 = data_d1[143:136];
        5'd19: vec_data_024 = data_d1[151:144];
        5'd20: vec_data_024 = data_d1[159:152];
        5'd21: vec_data_024 = data_d1[167:160];
        5'd22: vec_data_024 = data_d1[175:168];
        5'd23: vec_data_024 = data_d1[183:176];
        5'd24: vec_data_024 = data_d1[191:184];
        5'd25: vec_data_024 = data_d1[199:192];
    endcase
end

always @(
  vec_sum_025_d1
  or data_d1
  ) begin
    vec_data_025 = 8'b0;
    case(vec_sum_025_d1)
        5'd1: vec_data_025 = data_d1[7:0];
        5'd2: vec_data_025 = data_d1[15:8];
        5'd3: vec_data_025 = data_d1[23:16];
        5'd4: vec_data_025 = data_d1[31:24];
        5'd5: vec_data_025 = data_d1[39:32];
        5'd6: vec_data_025 = data_d1[47:40];
        5'd7: vec_data_025 = data_d1[55:48];
        5'd8: vec_data_025 = data_d1[63:56];
        5'd9: vec_data_025 = data_d1[71:64];
        5'd10: vec_data_025 = data_d1[79:72];
        5'd11: vec_data_025 = data_d1[87:80];
        5'd12: vec_data_025 = data_d1[95:88];
        5'd13: vec_data_025 = data_d1[103:96];
        5'd14: vec_data_025 = data_d1[111:104];
        5'd15: vec_data_025 = data_d1[119:112];
        5'd16: vec_data_025 = data_d1[127:120];
        5'd17: vec_data_025 = data_d1[135:128];
        5'd18: vec_data_025 = data_d1[143:136];
        5'd19: vec_data_025 = data_d1[151:144];
        5'd20: vec_data_025 = data_d1[159:152];
        5'd21: vec_data_025 = data_d1[167:160];
        5'd22: vec_data_025 = data_d1[175:168];
        5'd23: vec_data_025 = data_d1[183:176];
        5'd24: vec_data_025 = data_d1[191:184];
        5'd25: vec_data_025 = data_d1[199:192];
        5'd26: vec_data_025 = data_d1[207:200];
    endcase
end

always @(
  vec_sum_026_d1
  or data_d1
  ) begin
    vec_data_026 = 8'b0;
    case(vec_sum_026_d1)
        5'd1: vec_data_026 = data_d1[7:0];
        5'd2: vec_data_026 = data_d1[15:8];
        5'd3: vec_data_026 = data_d1[23:16];
        5'd4: vec_data_026 = data_d1[31:24];
        5'd5: vec_data_026 = data_d1[39:32];
        5'd6: vec_data_026 = data_d1[47:40];
        5'd7: vec_data_026 = data_d1[55:48];
        5'd8: vec_data_026 = data_d1[63:56];
        5'd9: vec_data_026 = data_d1[71:64];
        5'd10: vec_data_026 = data_d1[79:72];
        5'd11: vec_data_026 = data_d1[87:80];
        5'd12: vec_data_026 = data_d1[95:88];
        5'd13: vec_data_026 = data_d1[103:96];
        5'd14: vec_data_026 = data_d1[111:104];
        5'd15: vec_data_026 = data_d1[119:112];
        5'd16: vec_data_026 = data_d1[127:120];
        5'd17: vec_data_026 = data_d1[135:128];
        5'd18: vec_data_026 = data_d1[143:136];
        5'd19: vec_data_026 = data_d1[151:144];
        5'd20: vec_data_026 = data_d1[159:152];
        5'd21: vec_data_026 = data_d1[167:160];
        5'd22: vec_data_026 = data_d1[175:168];
        5'd23: vec_data_026 = data_d1[183:176];
        5'd24: vec_data_026 = data_d1[191:184];
        5'd25: vec_data_026 = data_d1[199:192];
        5'd26: vec_data_026 = data_d1[207:200];
        5'd27: vec_data_026 = data_d1[215:208];
    endcase
end

always @(
  vec_sum_027_d1
  or data_d1
  ) begin
    vec_data_027 = 8'b0;
    case(vec_sum_027_d1)
        5'd1: vec_data_027 = data_d1[7:0];
        5'd2: vec_data_027 = data_d1[15:8];
        5'd3: vec_data_027 = data_d1[23:16];
        5'd4: vec_data_027 = data_d1[31:24];
        5'd5: vec_data_027 = data_d1[39:32];
        5'd6: vec_data_027 = data_d1[47:40];
        5'd7: vec_data_027 = data_d1[55:48];
        5'd8: vec_data_027 = data_d1[63:56];
        5'd9: vec_data_027 = data_d1[71:64];
        5'd10: vec_data_027 = data_d1[79:72];
        5'd11: vec_data_027 = data_d1[87:80];
        5'd12: vec_data_027 = data_d1[95:88];
        5'd13: vec_data_027 = data_d1[103:96];
        5'd14: vec_data_027 = data_d1[111:104];
        5'd15: vec_data_027 = data_d1[119:112];
        5'd16: vec_data_027 = data_d1[127:120];
        5'd17: vec_data_027 = data_d1[135:128];
        5'd18: vec_data_027 = data_d1[143:136];
        5'd19: vec_data_027 = data_d1[151:144];
        5'd20: vec_data_027 = data_d1[159:152];
        5'd21: vec_data_027 = data_d1[167:160];
        5'd22: vec_data_027 = data_d1[175:168];
        5'd23: vec_data_027 = data_d1[183:176];
        5'd24: vec_data_027 = data_d1[191:184];
        5'd25: vec_data_027 = data_d1[199:192];
        5'd26: vec_data_027 = data_d1[207:200];
        5'd27: vec_data_027 = data_d1[215:208];
        5'd28: vec_data_027 = data_d1[223:216];
    endcase
end

always @(
  vec_sum_028_d1
  or data_d1
  ) begin
    vec_data_028 = 8'b0;
    case(vec_sum_028_d1)
        5'd1: vec_data_028 = data_d1[7:0];
        5'd2: vec_data_028 = data_d1[15:8];
        5'd3: vec_data_028 = data_d1[23:16];
        5'd4: vec_data_028 = data_d1[31:24];
        5'd5: vec_data_028 = data_d1[39:32];
        5'd6: vec_data_028 = data_d1[47:40];
        5'd7: vec_data_028 = data_d1[55:48];
        5'd8: vec_data_028 = data_d1[63:56];
        5'd9: vec_data_028 = data_d1[71:64];
        5'd10: vec_data_028 = data_d1[79:72];
        5'd11: vec_data_028 = data_d1[87:80];
        5'd12: vec_data_028 = data_d1[95:88];
        5'd13: vec_data_028 = data_d1[103:96];
        5'd14: vec_data_028 = data_d1[111:104];
        5'd15: vec_data_028 = data_d1[119:112];
        5'd16: vec_data_028 = data_d1[127:120];
        5'd17: vec_data_028 = data_d1[135:128];
        5'd18: vec_data_028 = data_d1[143:136];
        5'd19: vec_data_028 = data_d1[151:144];
        5'd20: vec_data_028 = data_d1[159:152];
        5'd21: vec_data_028 = data_d1[167:160];
        5'd22: vec_data_028 = data_d1[175:168];
        5'd23: vec_data_028 = data_d1[183:176];
        5'd24: vec_data_028 = data_d1[191:184];
        5'd25: vec_data_028 = data_d1[199:192];
        5'd26: vec_data_028 = data_d1[207:200];
        5'd27: vec_data_028 = data_d1[215:208];
        5'd28: vec_data_028 = data_d1[223:216];
        5'd29: vec_data_028 = data_d1[231:224];
    endcase
end

always @(
  vec_sum_029_d1
  or data_d1
  ) begin
    vec_data_029 = 8'b0;
    case(vec_sum_029_d1)
        5'd1: vec_data_029 = data_d1[7:0];
        5'd2: vec_data_029 = data_d1[15:8];
        5'd3: vec_data_029 = data_d1[23:16];
        5'd4: vec_data_029 = data_d1[31:24];
        5'd5: vec_data_029 = data_d1[39:32];
        5'd6: vec_data_029 = data_d1[47:40];
        5'd7: vec_data_029 = data_d1[55:48];
        5'd8: vec_data_029 = data_d1[63:56];
        5'd9: vec_data_029 = data_d1[71:64];
        5'd10: vec_data_029 = data_d1[79:72];
        5'd11: vec_data_029 = data_d1[87:80];
        5'd12: vec_data_029 = data_d1[95:88];
        5'd13: vec_data_029 = data_d1[103:96];
        5'd14: vec_data_029 = data_d1[111:104];
        5'd15: vec_data_029 = data_d1[119:112];
        5'd16: vec_data_029 = data_d1[127:120];
        5'd17: vec_data_029 = data_d1[135:128];
        5'd18: vec_data_029 = data_d1[143:136];
        5'd19: vec_data_029 = data_d1[151:144];
        5'd20: vec_data_029 = data_d1[159:152];
        5'd21: vec_data_029 = data_d1[167:160];
        5'd22: vec_data_029 = data_d1[175:168];
        5'd23: vec_data_029 = data_d1[183:176];
        5'd24: vec_data_029 = data_d1[191:184];
        5'd25: vec_data_029 = data_d1[199:192];
        5'd26: vec_data_029 = data_d1[207:200];
        5'd27: vec_data_029 = data_d1[215:208];
        5'd28: vec_data_029 = data_d1[223:216];
        5'd29: vec_data_029 = data_d1[231:224];
        5'd30: vec_data_029 = data_d1[239:232];
    endcase
end

always @(
  vec_sum_030_d1
  or data_d1
  ) begin
    vec_data_030 = 8'b0;
    case(vec_sum_030_d1)
        5'd1: vec_data_030 = data_d1[7:0];
        5'd2: vec_data_030 = data_d1[15:8];
        5'd3: vec_data_030 = data_d1[23:16];
        5'd4: vec_data_030 = data_d1[31:24];
        5'd5: vec_data_030 = data_d1[39:32];
        5'd6: vec_data_030 = data_d1[47:40];
        5'd7: vec_data_030 = data_d1[55:48];
        5'd8: vec_data_030 = data_d1[63:56];
        5'd9: vec_data_030 = data_d1[71:64];
        5'd10: vec_data_030 = data_d1[79:72];
        5'd11: vec_data_030 = data_d1[87:80];
        5'd12: vec_data_030 = data_d1[95:88];
        5'd13: vec_data_030 = data_d1[103:96];
        5'd14: vec_data_030 = data_d1[111:104];
        5'd15: vec_data_030 = data_d1[119:112];
        5'd16: vec_data_030 = data_d1[127:120];
        5'd17: vec_data_030 = data_d1[135:128];
        5'd18: vec_data_030 = data_d1[143:136];
        5'd19: vec_data_030 = data_d1[151:144];
        5'd20: vec_data_030 = data_d1[159:152];
        5'd21: vec_data_030 = data_d1[167:160];
        5'd22: vec_data_030 = data_d1[175:168];
        5'd23: vec_data_030 = data_d1[183:176];
        5'd24: vec_data_030 = data_d1[191:184];
        5'd25: vec_data_030 = data_d1[199:192];
        5'd26: vec_data_030 = data_d1[207:200];
        5'd27: vec_data_030 = data_d1[215:208];
        5'd28: vec_data_030 = data_d1[223:216];
        5'd29: vec_data_030 = data_d1[231:224];
        5'd30: vec_data_030 = data_d1[239:232];
        5'd31: vec_data_030 = data_d1[247:240];
    endcase
end

always @(
  vec_sum_031_d1
  or data_d1
  ) begin
    vec_data_031 = 8'b0;
    case(vec_sum_031_d1)
        6'd1: vec_data_031 = data_d1[7:0];
        6'd2: vec_data_031 = data_d1[15:8];
        6'd3: vec_data_031 = data_d1[23:16];
        6'd4: vec_data_031 = data_d1[31:24];
        6'd5: vec_data_031 = data_d1[39:32];
        6'd6: vec_data_031 = data_d1[47:40];
        6'd7: vec_data_031 = data_d1[55:48];
        6'd8: vec_data_031 = data_d1[63:56];
        6'd9: vec_data_031 = data_d1[71:64];
        6'd10: vec_data_031 = data_d1[79:72];
        6'd11: vec_data_031 = data_d1[87:80];
        6'd12: vec_data_031 = data_d1[95:88];
        6'd13: vec_data_031 = data_d1[103:96];
        6'd14: vec_data_031 = data_d1[111:104];
        6'd15: vec_data_031 = data_d1[119:112];
        6'd16: vec_data_031 = data_d1[127:120];
        6'd17: vec_data_031 = data_d1[135:128];
        6'd18: vec_data_031 = data_d1[143:136];
        6'd19: vec_data_031 = data_d1[151:144];
        6'd20: vec_data_031 = data_d1[159:152];
        6'd21: vec_data_031 = data_d1[167:160];
        6'd22: vec_data_031 = data_d1[175:168];
        6'd23: vec_data_031 = data_d1[183:176];
        6'd24: vec_data_031 = data_d1[191:184];
        6'd25: vec_data_031 = data_d1[199:192];
        6'd26: vec_data_031 = data_d1[207:200];
        6'd27: vec_data_031 = data_d1[215:208];
        6'd28: vec_data_031 = data_d1[223:216];
        6'd29: vec_data_031 = data_d1[231:224];
        6'd30: vec_data_031 = data_d1[239:232];
        6'd31: vec_data_031 = data_d1[247:240];
        6'd32: vec_data_031 = data_d1[255:248];
    endcase
end

always @(
  vec_sum_032_d1
  or data_d1
  ) begin
    vec_data_032 = 8'b0;
    case(vec_sum_032_d1)
        6'd1: vec_data_032 = data_d1[7:0];
        6'd2: vec_data_032 = data_d1[15:8];
        6'd3: vec_data_032 = data_d1[23:16];
        6'd4: vec_data_032 = data_d1[31:24];
        6'd5: vec_data_032 = data_d1[39:32];
        6'd6: vec_data_032 = data_d1[47:40];
        6'd7: vec_data_032 = data_d1[55:48];
        6'd8: vec_data_032 = data_d1[63:56];
        6'd9: vec_data_032 = data_d1[71:64];
        6'd10: vec_data_032 = data_d1[79:72];
        6'd11: vec_data_032 = data_d1[87:80];
        6'd12: vec_data_032 = data_d1[95:88];
        6'd13: vec_data_032 = data_d1[103:96];
        6'd14: vec_data_032 = data_d1[111:104];
        6'd15: vec_data_032 = data_d1[119:112];
        6'd16: vec_data_032 = data_d1[127:120];
        6'd17: vec_data_032 = data_d1[135:128];
        6'd18: vec_data_032 = data_d1[143:136];
        6'd19: vec_data_032 = data_d1[151:144];
        6'd20: vec_data_032 = data_d1[159:152];
        6'd21: vec_data_032 = data_d1[167:160];
        6'd22: vec_data_032 = data_d1[175:168];
        6'd23: vec_data_032 = data_d1[183:176];
        6'd24: vec_data_032 = data_d1[191:184];
        6'd25: vec_data_032 = data_d1[199:192];
        6'd26: vec_data_032 = data_d1[207:200];
        6'd27: vec_data_032 = data_d1[215:208];
        6'd28: vec_data_032 = data_d1[223:216];
        6'd29: vec_data_032 = data_d1[231:224];
        6'd30: vec_data_032 = data_d1[239:232];
        6'd31: vec_data_032 = data_d1[247:240];
        6'd32: vec_data_032 = data_d1[255:248];
        6'd33: vec_data_032 = data_d1[263:256];
    endcase
end

always @(
  vec_sum_033_d1
  or data_d1
  ) begin
    vec_data_033 = 8'b0;
    case(vec_sum_033_d1)
        6'd1: vec_data_033 = data_d1[7:0];
        6'd2: vec_data_033 = data_d1[15:8];
        6'd3: vec_data_033 = data_d1[23:16];
        6'd4: vec_data_033 = data_d1[31:24];
        6'd5: vec_data_033 = data_d1[39:32];
        6'd6: vec_data_033 = data_d1[47:40];
        6'd7: vec_data_033 = data_d1[55:48];
        6'd8: vec_data_033 = data_d1[63:56];
        6'd9: vec_data_033 = data_d1[71:64];
        6'd10: vec_data_033 = data_d1[79:72];
        6'd11: vec_data_033 = data_d1[87:80];
        6'd12: vec_data_033 = data_d1[95:88];
        6'd13: vec_data_033 = data_d1[103:96];
        6'd14: vec_data_033 = data_d1[111:104];
        6'd15: vec_data_033 = data_d1[119:112];
        6'd16: vec_data_033 = data_d1[127:120];
        6'd17: vec_data_033 = data_d1[135:128];
        6'd18: vec_data_033 = data_d1[143:136];
        6'd19: vec_data_033 = data_d1[151:144];
        6'd20: vec_data_033 = data_d1[159:152];
        6'd21: vec_data_033 = data_d1[167:160];
        6'd22: vec_data_033 = data_d1[175:168];
        6'd23: vec_data_033 = data_d1[183:176];
        6'd24: vec_data_033 = data_d1[191:184];
        6'd25: vec_data_033 = data_d1[199:192];
        6'd26: vec_data_033 = data_d1[207:200];
        6'd27: vec_data_033 = data_d1[215:208];
        6'd28: vec_data_033 = data_d1[223:216];
        6'd29: vec_data_033 = data_d1[231:224];
        6'd30: vec_data_033 = data_d1[239:232];
        6'd31: vec_data_033 = data_d1[247:240];
        6'd32: vec_data_033 = data_d1[255:248];
        6'd33: vec_data_033 = data_d1[263:256];
        6'd34: vec_data_033 = data_d1[271:264];
    endcase
end

always @(
  vec_sum_034_d1
  or data_d1
  ) begin
    vec_data_034 = 8'b0;
    case(vec_sum_034_d1)
        6'd1: vec_data_034 = data_d1[7:0];
        6'd2: vec_data_034 = data_d1[15:8];
        6'd3: vec_data_034 = data_d1[23:16];
        6'd4: vec_data_034 = data_d1[31:24];
        6'd5: vec_data_034 = data_d1[39:32];
        6'd6: vec_data_034 = data_d1[47:40];
        6'd7: vec_data_034 = data_d1[55:48];
        6'd8: vec_data_034 = data_d1[63:56];
        6'd9: vec_data_034 = data_d1[71:64];
        6'd10: vec_data_034 = data_d1[79:72];
        6'd11: vec_data_034 = data_d1[87:80];
        6'd12: vec_data_034 = data_d1[95:88];
        6'd13: vec_data_034 = data_d1[103:96];
        6'd14: vec_data_034 = data_d1[111:104];
        6'd15: vec_data_034 = data_d1[119:112];
        6'd16: vec_data_034 = data_d1[127:120];
        6'd17: vec_data_034 = data_d1[135:128];
        6'd18: vec_data_034 = data_d1[143:136];
        6'd19: vec_data_034 = data_d1[151:144];
        6'd20: vec_data_034 = data_d1[159:152];
        6'd21: vec_data_034 = data_d1[167:160];
        6'd22: vec_data_034 = data_d1[175:168];
        6'd23: vec_data_034 = data_d1[183:176];
        6'd24: vec_data_034 = data_d1[191:184];
        6'd25: vec_data_034 = data_d1[199:192];
        6'd26: vec_data_034 = data_d1[207:200];
        6'd27: vec_data_034 = data_d1[215:208];
        6'd28: vec_data_034 = data_d1[223:216];
        6'd29: vec_data_034 = data_d1[231:224];
        6'd30: vec_data_034 = data_d1[239:232];
        6'd31: vec_data_034 = data_d1[247:240];
        6'd32: vec_data_034 = data_d1[255:248];
        6'd33: vec_data_034 = data_d1[263:256];
        6'd34: vec_data_034 = data_d1[271:264];
        6'd35: vec_data_034 = data_d1[279:272];
    endcase
end

always @(
  vec_sum_035_d1
  or data_d1
  ) begin
    vec_data_035 = 8'b0;
    case(vec_sum_035_d1)
        6'd1: vec_data_035 = data_d1[7:0];
        6'd2: vec_data_035 = data_d1[15:8];
        6'd3: vec_data_035 = data_d1[23:16];
        6'd4: vec_data_035 = data_d1[31:24];
        6'd5: vec_data_035 = data_d1[39:32];
        6'd6: vec_data_035 = data_d1[47:40];
        6'd7: vec_data_035 = data_d1[55:48];
        6'd8: vec_data_035 = data_d1[63:56];
        6'd9: vec_data_035 = data_d1[71:64];
        6'd10: vec_data_035 = data_d1[79:72];
        6'd11: vec_data_035 = data_d1[87:80];
        6'd12: vec_data_035 = data_d1[95:88];
        6'd13: vec_data_035 = data_d1[103:96];
        6'd14: vec_data_035 = data_d1[111:104];
        6'd15: vec_data_035 = data_d1[119:112];
        6'd16: vec_data_035 = data_d1[127:120];
        6'd17: vec_data_035 = data_d1[135:128];
        6'd18: vec_data_035 = data_d1[143:136];
        6'd19: vec_data_035 = data_d1[151:144];
        6'd20: vec_data_035 = data_d1[159:152];
        6'd21: vec_data_035 = data_d1[167:160];
        6'd22: vec_data_035 = data_d1[175:168];
        6'd23: vec_data_035 = data_d1[183:176];
        6'd24: vec_data_035 = data_d1[191:184];
        6'd25: vec_data_035 = data_d1[199:192];
        6'd26: vec_data_035 = data_d1[207:200];
        6'd27: vec_data_035 = data_d1[215:208];
        6'd28: vec_data_035 = data_d1[223:216];
        6'd29: vec_data_035 = data_d1[231:224];
        6'd30: vec_data_035 = data_d1[239:232];
        6'd31: vec_data_035 = data_d1[247:240];
        6'd32: vec_data_035 = data_d1[255:248];
        6'd33: vec_data_035 = data_d1[263:256];
        6'd34: vec_data_035 = data_d1[271:264];
        6'd35: vec_data_035 = data_d1[279:272];
        6'd36: vec_data_035 = data_d1[287:280];
    endcase
end

always @(
  vec_sum_036_d1
  or data_d1
  ) begin
    vec_data_036 = 8'b0;
    case(vec_sum_036_d1)
        6'd1: vec_data_036 = data_d1[7:0];
        6'd2: vec_data_036 = data_d1[15:8];
        6'd3: vec_data_036 = data_d1[23:16];
        6'd4: vec_data_036 = data_d1[31:24];
        6'd5: vec_data_036 = data_d1[39:32];
        6'd6: vec_data_036 = data_d1[47:40];
        6'd7: vec_data_036 = data_d1[55:48];
        6'd8: vec_data_036 = data_d1[63:56];
        6'd9: vec_data_036 = data_d1[71:64];
        6'd10: vec_data_036 = data_d1[79:72];
        6'd11: vec_data_036 = data_d1[87:80];
        6'd12: vec_data_036 = data_d1[95:88];
        6'd13: vec_data_036 = data_d1[103:96];
        6'd14: vec_data_036 = data_d1[111:104];
        6'd15: vec_data_036 = data_d1[119:112];
        6'd16: vec_data_036 = data_d1[127:120];
        6'd17: vec_data_036 = data_d1[135:128];
        6'd18: vec_data_036 = data_d1[143:136];
        6'd19: vec_data_036 = data_d1[151:144];
        6'd20: vec_data_036 = data_d1[159:152];
        6'd21: vec_data_036 = data_d1[167:160];
        6'd22: vec_data_036 = data_d1[175:168];
        6'd23: vec_data_036 = data_d1[183:176];
        6'd24: vec_data_036 = data_d1[191:184];
        6'd25: vec_data_036 = data_d1[199:192];
        6'd26: vec_data_036 = data_d1[207:200];
        6'd27: vec_data_036 = data_d1[215:208];
        6'd28: vec_data_036 = data_d1[223:216];
        6'd29: vec_data_036 = data_d1[231:224];
        6'd30: vec_data_036 = data_d1[239:232];
        6'd31: vec_data_036 = data_d1[247:240];
        6'd32: vec_data_036 = data_d1[255:248];
        6'd33: vec_data_036 = data_d1[263:256];
        6'd34: vec_data_036 = data_d1[271:264];
        6'd35: vec_data_036 = data_d1[279:272];
        6'd36: vec_data_036 = data_d1[287:280];
        6'd37: vec_data_036 = data_d1[295:288];
    endcase
end

always @(
  vec_sum_037_d1
  or data_d1
  ) begin
    vec_data_037 = 8'b0;
    case(vec_sum_037_d1)
        6'd1: vec_data_037 = data_d1[7:0];
        6'd2: vec_data_037 = data_d1[15:8];
        6'd3: vec_data_037 = data_d1[23:16];
        6'd4: vec_data_037 = data_d1[31:24];
        6'd5: vec_data_037 = data_d1[39:32];
        6'd6: vec_data_037 = data_d1[47:40];
        6'd7: vec_data_037 = data_d1[55:48];
        6'd8: vec_data_037 = data_d1[63:56];
        6'd9: vec_data_037 = data_d1[71:64];
        6'd10: vec_data_037 = data_d1[79:72];
        6'd11: vec_data_037 = data_d1[87:80];
        6'd12: vec_data_037 = data_d1[95:88];
        6'd13: vec_data_037 = data_d1[103:96];
        6'd14: vec_data_037 = data_d1[111:104];
        6'd15: vec_data_037 = data_d1[119:112];
        6'd16: vec_data_037 = data_d1[127:120];
        6'd17: vec_data_037 = data_d1[135:128];
        6'd18: vec_data_037 = data_d1[143:136];
        6'd19: vec_data_037 = data_d1[151:144];
        6'd20: vec_data_037 = data_d1[159:152];
        6'd21: vec_data_037 = data_d1[167:160];
        6'd22: vec_data_037 = data_d1[175:168];
        6'd23: vec_data_037 = data_d1[183:176];
        6'd24: vec_data_037 = data_d1[191:184];
        6'd25: vec_data_037 = data_d1[199:192];
        6'd26: vec_data_037 = data_d1[207:200];
        6'd27: vec_data_037 = data_d1[215:208];
        6'd28: vec_data_037 = data_d1[223:216];
        6'd29: vec_data_037 = data_d1[231:224];
        6'd30: vec_data_037 = data_d1[239:232];
        6'd31: vec_data_037 = data_d1[247:240];
        6'd32: vec_data_037 = data_d1[255:248];
        6'd33: vec_data_037 = data_d1[263:256];
        6'd34: vec_data_037 = data_d1[271:264];
        6'd35: vec_data_037 = data_d1[279:272];
        6'd36: vec_data_037 = data_d1[287:280];
        6'd37: vec_data_037 = data_d1[295:288];
        6'd38: vec_data_037 = data_d1[303:296];
    endcase
end

always @(
  vec_sum_038_d1
  or data_d1
  ) begin
    vec_data_038 = 8'b0;
    case(vec_sum_038_d1)
        6'd1: vec_data_038 = data_d1[7:0];
        6'd2: vec_data_038 = data_d1[15:8];
        6'd3: vec_data_038 = data_d1[23:16];
        6'd4: vec_data_038 = data_d1[31:24];
        6'd5: vec_data_038 = data_d1[39:32];
        6'd6: vec_data_038 = data_d1[47:40];
        6'd7: vec_data_038 = data_d1[55:48];
        6'd8: vec_data_038 = data_d1[63:56];
        6'd9: vec_data_038 = data_d1[71:64];
        6'd10: vec_data_038 = data_d1[79:72];
        6'd11: vec_data_038 = data_d1[87:80];
        6'd12: vec_data_038 = data_d1[95:88];
        6'd13: vec_data_038 = data_d1[103:96];
        6'd14: vec_data_038 = data_d1[111:104];
        6'd15: vec_data_038 = data_d1[119:112];
        6'd16: vec_data_038 = data_d1[127:120];
        6'd17: vec_data_038 = data_d1[135:128];
        6'd18: vec_data_038 = data_d1[143:136];
        6'd19: vec_data_038 = data_d1[151:144];
        6'd20: vec_data_038 = data_d1[159:152];
        6'd21: vec_data_038 = data_d1[167:160];
        6'd22: vec_data_038 = data_d1[175:168];
        6'd23: vec_data_038 = data_d1[183:176];
        6'd24: vec_data_038 = data_d1[191:184];
        6'd25: vec_data_038 = data_d1[199:192];
        6'd26: vec_data_038 = data_d1[207:200];
        6'd27: vec_data_038 = data_d1[215:208];
        6'd28: vec_data_038 = data_d1[223:216];
        6'd29: vec_data_038 = data_d1[231:224];
        6'd30: vec_data_038 = data_d1[239:232];
        6'd31: vec_data_038 = data_d1[247:240];
        6'd32: vec_data_038 = data_d1[255:248];
        6'd33: vec_data_038 = data_d1[263:256];
        6'd34: vec_data_038 = data_d1[271:264];
        6'd35: vec_data_038 = data_d1[279:272];
        6'd36: vec_data_038 = data_d1[287:280];
        6'd37: vec_data_038 = data_d1[295:288];
        6'd38: vec_data_038 = data_d1[303:296];
        6'd39: vec_data_038 = data_d1[311:304];
    endcase
end

always @(
  vec_sum_039_d1
  or data_d1
  ) begin
    vec_data_039 = 8'b0;
    case(vec_sum_039_d1)
        6'd1: vec_data_039 = data_d1[7:0];
        6'd2: vec_data_039 = data_d1[15:8];
        6'd3: vec_data_039 = data_d1[23:16];
        6'd4: vec_data_039 = data_d1[31:24];
        6'd5: vec_data_039 = data_d1[39:32];
        6'd6: vec_data_039 = data_d1[47:40];
        6'd7: vec_data_039 = data_d1[55:48];
        6'd8: vec_data_039 = data_d1[63:56];
        6'd9: vec_data_039 = data_d1[71:64];
        6'd10: vec_data_039 = data_d1[79:72];
        6'd11: vec_data_039 = data_d1[87:80];
        6'd12: vec_data_039 = data_d1[95:88];
        6'd13: vec_data_039 = data_d1[103:96];
        6'd14: vec_data_039 = data_d1[111:104];
        6'd15: vec_data_039 = data_d1[119:112];
        6'd16: vec_data_039 = data_d1[127:120];
        6'd17: vec_data_039 = data_d1[135:128];
        6'd18: vec_data_039 = data_d1[143:136];
        6'd19: vec_data_039 = data_d1[151:144];
        6'd20: vec_data_039 = data_d1[159:152];
        6'd21: vec_data_039 = data_d1[167:160];
        6'd22: vec_data_039 = data_d1[175:168];
        6'd23: vec_data_039 = data_d1[183:176];
        6'd24: vec_data_039 = data_d1[191:184];
        6'd25: vec_data_039 = data_d1[199:192];
        6'd26: vec_data_039 = data_d1[207:200];
        6'd27: vec_data_039 = data_d1[215:208];
        6'd28: vec_data_039 = data_d1[223:216];
        6'd29: vec_data_039 = data_d1[231:224];
        6'd30: vec_data_039 = data_d1[239:232];
        6'd31: vec_data_039 = data_d1[247:240];
        6'd32: vec_data_039 = data_d1[255:248];
        6'd33: vec_data_039 = data_d1[263:256];
        6'd34: vec_data_039 = data_d1[271:264];
        6'd35: vec_data_039 = data_d1[279:272];
        6'd36: vec_data_039 = data_d1[287:280];
        6'd37: vec_data_039 = data_d1[295:288];
        6'd38: vec_data_039 = data_d1[303:296];
        6'd39: vec_data_039 = data_d1[311:304];
        6'd40: vec_data_039 = data_d1[319:312];
    endcase
end

always @(
  vec_sum_040_d1
  or data_d1
  ) begin
    vec_data_040 = 8'b0;
    case(vec_sum_040_d1)
        6'd1: vec_data_040 = data_d1[7:0];
        6'd2: vec_data_040 = data_d1[15:8];
        6'd3: vec_data_040 = data_d1[23:16];
        6'd4: vec_data_040 = data_d1[31:24];
        6'd5: vec_data_040 = data_d1[39:32];
        6'd6: vec_data_040 = data_d1[47:40];
        6'd7: vec_data_040 = data_d1[55:48];
        6'd8: vec_data_040 = data_d1[63:56];
        6'd9: vec_data_040 = data_d1[71:64];
        6'd10: vec_data_040 = data_d1[79:72];
        6'd11: vec_data_040 = data_d1[87:80];
        6'd12: vec_data_040 = data_d1[95:88];
        6'd13: vec_data_040 = data_d1[103:96];
        6'd14: vec_data_040 = data_d1[111:104];
        6'd15: vec_data_040 = data_d1[119:112];
        6'd16: vec_data_040 = data_d1[127:120];
        6'd17: vec_data_040 = data_d1[135:128];
        6'd18: vec_data_040 = data_d1[143:136];
        6'd19: vec_data_040 = data_d1[151:144];
        6'd20: vec_data_040 = data_d1[159:152];
        6'd21: vec_data_040 = data_d1[167:160];
        6'd22: vec_data_040 = data_d1[175:168];
        6'd23: vec_data_040 = data_d1[183:176];
        6'd24: vec_data_040 = data_d1[191:184];
        6'd25: vec_data_040 = data_d1[199:192];
        6'd26: vec_data_040 = data_d1[207:200];
        6'd27: vec_data_040 = data_d1[215:208];
        6'd28: vec_data_040 = data_d1[223:216];
        6'd29: vec_data_040 = data_d1[231:224];
        6'd30: vec_data_040 = data_d1[239:232];
        6'd31: vec_data_040 = data_d1[247:240];
        6'd32: vec_data_040 = data_d1[255:248];
        6'd33: vec_data_040 = data_d1[263:256];
        6'd34: vec_data_040 = data_d1[271:264];
        6'd35: vec_data_040 = data_d1[279:272];
        6'd36: vec_data_040 = data_d1[287:280];
        6'd37: vec_data_040 = data_d1[295:288];
        6'd38: vec_data_040 = data_d1[303:296];
        6'd39: vec_data_040 = data_d1[311:304];
        6'd40: vec_data_040 = data_d1[319:312];
        6'd41: vec_data_040 = data_d1[327:320];
    endcase
end

always @(
  vec_sum_041_d1
  or data_d1
  ) begin
    vec_data_041 = 8'b0;
    case(vec_sum_041_d1)
        6'd1: vec_data_041 = data_d1[7:0];
        6'd2: vec_data_041 = data_d1[15:8];
        6'd3: vec_data_041 = data_d1[23:16];
        6'd4: vec_data_041 = data_d1[31:24];
        6'd5: vec_data_041 = data_d1[39:32];
        6'd6: vec_data_041 = data_d1[47:40];
        6'd7: vec_data_041 = data_d1[55:48];
        6'd8: vec_data_041 = data_d1[63:56];
        6'd9: vec_data_041 = data_d1[71:64];
        6'd10: vec_data_041 = data_d1[79:72];
        6'd11: vec_data_041 = data_d1[87:80];
        6'd12: vec_data_041 = data_d1[95:88];
        6'd13: vec_data_041 = data_d1[103:96];
        6'd14: vec_data_041 = data_d1[111:104];
        6'd15: vec_data_041 = data_d1[119:112];
        6'd16: vec_data_041 = data_d1[127:120];
        6'd17: vec_data_041 = data_d1[135:128];
        6'd18: vec_data_041 = data_d1[143:136];
        6'd19: vec_data_041 = data_d1[151:144];
        6'd20: vec_data_041 = data_d1[159:152];
        6'd21: vec_data_041 = data_d1[167:160];
        6'd22: vec_data_041 = data_d1[175:168];
        6'd23: vec_data_041 = data_d1[183:176];
        6'd24: vec_data_041 = data_d1[191:184];
        6'd25: vec_data_041 = data_d1[199:192];
        6'd26: vec_data_041 = data_d1[207:200];
        6'd27: vec_data_041 = data_d1[215:208];
        6'd28: vec_data_041 = data_d1[223:216];
        6'd29: vec_data_041 = data_d1[231:224];
        6'd30: vec_data_041 = data_d1[239:232];
        6'd31: vec_data_041 = data_d1[247:240];
        6'd32: vec_data_041 = data_d1[255:248];
        6'd33: vec_data_041 = data_d1[263:256];
        6'd34: vec_data_041 = data_d1[271:264];
        6'd35: vec_data_041 = data_d1[279:272];
        6'd36: vec_data_041 = data_d1[287:280];
        6'd37: vec_data_041 = data_d1[295:288];
        6'd38: vec_data_041 = data_d1[303:296];
        6'd39: vec_data_041 = data_d1[311:304];
        6'd40: vec_data_041 = data_d1[319:312];
        6'd41: vec_data_041 = data_d1[327:320];
        6'd42: vec_data_041 = data_d1[335:328];
    endcase
end

always @(
  vec_sum_042_d1
  or data_d1
  ) begin
    vec_data_042 = 8'b0;
    case(vec_sum_042_d1)
        6'd1: vec_data_042 = data_d1[7:0];
        6'd2: vec_data_042 = data_d1[15:8];
        6'd3: vec_data_042 = data_d1[23:16];
        6'd4: vec_data_042 = data_d1[31:24];
        6'd5: vec_data_042 = data_d1[39:32];
        6'd6: vec_data_042 = data_d1[47:40];
        6'd7: vec_data_042 = data_d1[55:48];
        6'd8: vec_data_042 = data_d1[63:56];
        6'd9: vec_data_042 = data_d1[71:64];
        6'd10: vec_data_042 = data_d1[79:72];
        6'd11: vec_data_042 = data_d1[87:80];
        6'd12: vec_data_042 = data_d1[95:88];
        6'd13: vec_data_042 = data_d1[103:96];
        6'd14: vec_data_042 = data_d1[111:104];
        6'd15: vec_data_042 = data_d1[119:112];
        6'd16: vec_data_042 = data_d1[127:120];
        6'd17: vec_data_042 = data_d1[135:128];
        6'd18: vec_data_042 = data_d1[143:136];
        6'd19: vec_data_042 = data_d1[151:144];
        6'd20: vec_data_042 = data_d1[159:152];
        6'd21: vec_data_042 = data_d1[167:160];
        6'd22: vec_data_042 = data_d1[175:168];
        6'd23: vec_data_042 = data_d1[183:176];
        6'd24: vec_data_042 = data_d1[191:184];
        6'd25: vec_data_042 = data_d1[199:192];
        6'd26: vec_data_042 = data_d1[207:200];
        6'd27: vec_data_042 = data_d1[215:208];
        6'd28: vec_data_042 = data_d1[223:216];
        6'd29: vec_data_042 = data_d1[231:224];
        6'd30: vec_data_042 = data_d1[239:232];
        6'd31: vec_data_042 = data_d1[247:240];
        6'd32: vec_data_042 = data_d1[255:248];
        6'd33: vec_data_042 = data_d1[263:256];
        6'd34: vec_data_042 = data_d1[271:264];
        6'd35: vec_data_042 = data_d1[279:272];
        6'd36: vec_data_042 = data_d1[287:280];
        6'd37: vec_data_042 = data_d1[295:288];
        6'd38: vec_data_042 = data_d1[303:296];
        6'd39: vec_data_042 = data_d1[311:304];
        6'd40: vec_data_042 = data_d1[319:312];
        6'd41: vec_data_042 = data_d1[327:320];
        6'd42: vec_data_042 = data_d1[335:328];
        6'd43: vec_data_042 = data_d1[343:336];
    endcase
end

always @(
  vec_sum_043_d1
  or data_d1
  ) begin
    vec_data_043 = 8'b0;
    case(vec_sum_043_d1)
        6'd1: vec_data_043 = data_d1[7:0];
        6'd2: vec_data_043 = data_d1[15:8];
        6'd3: vec_data_043 = data_d1[23:16];
        6'd4: vec_data_043 = data_d1[31:24];
        6'd5: vec_data_043 = data_d1[39:32];
        6'd6: vec_data_043 = data_d1[47:40];
        6'd7: vec_data_043 = data_d1[55:48];
        6'd8: vec_data_043 = data_d1[63:56];
        6'd9: vec_data_043 = data_d1[71:64];
        6'd10: vec_data_043 = data_d1[79:72];
        6'd11: vec_data_043 = data_d1[87:80];
        6'd12: vec_data_043 = data_d1[95:88];
        6'd13: vec_data_043 = data_d1[103:96];
        6'd14: vec_data_043 = data_d1[111:104];
        6'd15: vec_data_043 = data_d1[119:112];
        6'd16: vec_data_043 = data_d1[127:120];
        6'd17: vec_data_043 = data_d1[135:128];
        6'd18: vec_data_043 = data_d1[143:136];
        6'd19: vec_data_043 = data_d1[151:144];
        6'd20: vec_data_043 = data_d1[159:152];
        6'd21: vec_data_043 = data_d1[167:160];
        6'd22: vec_data_043 = data_d1[175:168];
        6'd23: vec_data_043 = data_d1[183:176];
        6'd24: vec_data_043 = data_d1[191:184];
        6'd25: vec_data_043 = data_d1[199:192];
        6'd26: vec_data_043 = data_d1[207:200];
        6'd27: vec_data_043 = data_d1[215:208];
        6'd28: vec_data_043 = data_d1[223:216];
        6'd29: vec_data_043 = data_d1[231:224];
        6'd30: vec_data_043 = data_d1[239:232];
        6'd31: vec_data_043 = data_d1[247:240];
        6'd32: vec_data_043 = data_d1[255:248];
        6'd33: vec_data_043 = data_d1[263:256];
        6'd34: vec_data_043 = data_d1[271:264];
        6'd35: vec_data_043 = data_d1[279:272];
        6'd36: vec_data_043 = data_d1[287:280];
        6'd37: vec_data_043 = data_d1[295:288];
        6'd38: vec_data_043 = data_d1[303:296];
        6'd39: vec_data_043 = data_d1[311:304];
        6'd40: vec_data_043 = data_d1[319:312];
        6'd41: vec_data_043 = data_d1[327:320];
        6'd42: vec_data_043 = data_d1[335:328];
        6'd43: vec_data_043 = data_d1[343:336];
        6'd44: vec_data_043 = data_d1[351:344];
    endcase
end

always @(
  vec_sum_044_d1
  or data_d1
  ) begin
    vec_data_044 = 8'b0;
    case(vec_sum_044_d1)
        6'd1: vec_data_044 = data_d1[7:0];
        6'd2: vec_data_044 = data_d1[15:8];
        6'd3: vec_data_044 = data_d1[23:16];
        6'd4: vec_data_044 = data_d1[31:24];
        6'd5: vec_data_044 = data_d1[39:32];
        6'd6: vec_data_044 = data_d1[47:40];
        6'd7: vec_data_044 = data_d1[55:48];
        6'd8: vec_data_044 = data_d1[63:56];
        6'd9: vec_data_044 = data_d1[71:64];
        6'd10: vec_data_044 = data_d1[79:72];
        6'd11: vec_data_044 = data_d1[87:80];
        6'd12: vec_data_044 = data_d1[95:88];
        6'd13: vec_data_044 = data_d1[103:96];
        6'd14: vec_data_044 = data_d1[111:104];
        6'd15: vec_data_044 = data_d1[119:112];
        6'd16: vec_data_044 = data_d1[127:120];
        6'd17: vec_data_044 = data_d1[135:128];
        6'd18: vec_data_044 = data_d1[143:136];
        6'd19: vec_data_044 = data_d1[151:144];
        6'd20: vec_data_044 = data_d1[159:152];
        6'd21: vec_data_044 = data_d1[167:160];
        6'd22: vec_data_044 = data_d1[175:168];
        6'd23: vec_data_044 = data_d1[183:176];
        6'd24: vec_data_044 = data_d1[191:184];
        6'd25: vec_data_044 = data_d1[199:192];
        6'd26: vec_data_044 = data_d1[207:200];
        6'd27: vec_data_044 = data_d1[215:208];
        6'd28: vec_data_044 = data_d1[223:216];
        6'd29: vec_data_044 = data_d1[231:224];
        6'd30: vec_data_044 = data_d1[239:232];
        6'd31: vec_data_044 = data_d1[247:240];
        6'd32: vec_data_044 = data_d1[255:248];
        6'd33: vec_data_044 = data_d1[263:256];
        6'd34: vec_data_044 = data_d1[271:264];
        6'd35: vec_data_044 = data_d1[279:272];
        6'd36: vec_data_044 = data_d1[287:280];
        6'd37: vec_data_044 = data_d1[295:288];
        6'd38: vec_data_044 = data_d1[303:296];
        6'd39: vec_data_044 = data_d1[311:304];
        6'd40: vec_data_044 = data_d1[319:312];
        6'd41: vec_data_044 = data_d1[327:320];
        6'd42: vec_data_044 = data_d1[335:328];
        6'd43: vec_data_044 = data_d1[343:336];
        6'd44: vec_data_044 = data_d1[351:344];
        6'd45: vec_data_044 = data_d1[359:352];
    endcase
end

always @(
  vec_sum_045_d1
  or data_d1
  ) begin
    vec_data_045 = 8'b0;
    case(vec_sum_045_d1)
        6'd1: vec_data_045 = data_d1[7:0];
        6'd2: vec_data_045 = data_d1[15:8];
        6'd3: vec_data_045 = data_d1[23:16];
        6'd4: vec_data_045 = data_d1[31:24];
        6'd5: vec_data_045 = data_d1[39:32];
        6'd6: vec_data_045 = data_d1[47:40];
        6'd7: vec_data_045 = data_d1[55:48];
        6'd8: vec_data_045 = data_d1[63:56];
        6'd9: vec_data_045 = data_d1[71:64];
        6'd10: vec_data_045 = data_d1[79:72];
        6'd11: vec_data_045 = data_d1[87:80];
        6'd12: vec_data_045 = data_d1[95:88];
        6'd13: vec_data_045 = data_d1[103:96];
        6'd14: vec_data_045 = data_d1[111:104];
        6'd15: vec_data_045 = data_d1[119:112];
        6'd16: vec_data_045 = data_d1[127:120];
        6'd17: vec_data_045 = data_d1[135:128];
        6'd18: vec_data_045 = data_d1[143:136];
        6'd19: vec_data_045 = data_d1[151:144];
        6'd20: vec_data_045 = data_d1[159:152];
        6'd21: vec_data_045 = data_d1[167:160];
        6'd22: vec_data_045 = data_d1[175:168];
        6'd23: vec_data_045 = data_d1[183:176];
        6'd24: vec_data_045 = data_d1[191:184];
        6'd25: vec_data_045 = data_d1[199:192];
        6'd26: vec_data_045 = data_d1[207:200];
        6'd27: vec_data_045 = data_d1[215:208];
        6'd28: vec_data_045 = data_d1[223:216];
        6'd29: vec_data_045 = data_d1[231:224];
        6'd30: vec_data_045 = data_d1[239:232];
        6'd31: vec_data_045 = data_d1[247:240];
        6'd32: vec_data_045 = data_d1[255:248];
        6'd33: vec_data_045 = data_d1[263:256];
        6'd34: vec_data_045 = data_d1[271:264];
        6'd35: vec_data_045 = data_d1[279:272];
        6'd36: vec_data_045 = data_d1[287:280];
        6'd37: vec_data_045 = data_d1[295:288];
        6'd38: vec_data_045 = data_d1[303:296];
        6'd39: vec_data_045 = data_d1[311:304];
        6'd40: vec_data_045 = data_d1[319:312];
        6'd41: vec_data_045 = data_d1[327:320];
        6'd42: vec_data_045 = data_d1[335:328];
        6'd43: vec_data_045 = data_d1[343:336];
        6'd44: vec_data_045 = data_d1[351:344];
        6'd45: vec_data_045 = data_d1[359:352];
        6'd46: vec_data_045 = data_d1[367:360];
    endcase
end

always @(
  vec_sum_046_d1
  or data_d1
  ) begin
    vec_data_046 = 8'b0;
    case(vec_sum_046_d1)
        6'd1: vec_data_046 = data_d1[7:0];
        6'd2: vec_data_046 = data_d1[15:8];
        6'd3: vec_data_046 = data_d1[23:16];
        6'd4: vec_data_046 = data_d1[31:24];
        6'd5: vec_data_046 = data_d1[39:32];
        6'd6: vec_data_046 = data_d1[47:40];
        6'd7: vec_data_046 = data_d1[55:48];
        6'd8: vec_data_046 = data_d1[63:56];
        6'd9: vec_data_046 = data_d1[71:64];
        6'd10: vec_data_046 = data_d1[79:72];
        6'd11: vec_data_046 = data_d1[87:80];
        6'd12: vec_data_046 = data_d1[95:88];
        6'd13: vec_data_046 = data_d1[103:96];
        6'd14: vec_data_046 = data_d1[111:104];
        6'd15: vec_data_046 = data_d1[119:112];
        6'd16: vec_data_046 = data_d1[127:120];
        6'd17: vec_data_046 = data_d1[135:128];
        6'd18: vec_data_046 = data_d1[143:136];
        6'd19: vec_data_046 = data_d1[151:144];
        6'd20: vec_data_046 = data_d1[159:152];
        6'd21: vec_data_046 = data_d1[167:160];
        6'd22: vec_data_046 = data_d1[175:168];
        6'd23: vec_data_046 = data_d1[183:176];
        6'd24: vec_data_046 = data_d1[191:184];
        6'd25: vec_data_046 = data_d1[199:192];
        6'd26: vec_data_046 = data_d1[207:200];
        6'd27: vec_data_046 = data_d1[215:208];
        6'd28: vec_data_046 = data_d1[223:216];
        6'd29: vec_data_046 = data_d1[231:224];
        6'd30: vec_data_046 = data_d1[239:232];
        6'd31: vec_data_046 = data_d1[247:240];
        6'd32: vec_data_046 = data_d1[255:248];
        6'd33: vec_data_046 = data_d1[263:256];
        6'd34: vec_data_046 = data_d1[271:264];
        6'd35: vec_data_046 = data_d1[279:272];
        6'd36: vec_data_046 = data_d1[287:280];
        6'd37: vec_data_046 = data_d1[295:288];
        6'd38: vec_data_046 = data_d1[303:296];
        6'd39: vec_data_046 = data_d1[311:304];
        6'd40: vec_data_046 = data_d1[319:312];
        6'd41: vec_data_046 = data_d1[327:320];
        6'd42: vec_data_046 = data_d1[335:328];
        6'd43: vec_data_046 = data_d1[343:336];
        6'd44: vec_data_046 = data_d1[351:344];
        6'd45: vec_data_046 = data_d1[359:352];
        6'd46: vec_data_046 = data_d1[367:360];
        6'd47: vec_data_046 = data_d1[375:368];
    endcase
end

always @(
  vec_sum_047_d1
  or data_d1
  ) begin
    vec_data_047 = 8'b0;
    case(vec_sum_047_d1)
        6'd1: vec_data_047 = data_d1[7:0];
        6'd2: vec_data_047 = data_d1[15:8];
        6'd3: vec_data_047 = data_d1[23:16];
        6'd4: vec_data_047 = data_d1[31:24];
        6'd5: vec_data_047 = data_d1[39:32];
        6'd6: vec_data_047 = data_d1[47:40];
        6'd7: vec_data_047 = data_d1[55:48];
        6'd8: vec_data_047 = data_d1[63:56];
        6'd9: vec_data_047 = data_d1[71:64];
        6'd10: vec_data_047 = data_d1[79:72];
        6'd11: vec_data_047 = data_d1[87:80];
        6'd12: vec_data_047 = data_d1[95:88];
        6'd13: vec_data_047 = data_d1[103:96];
        6'd14: vec_data_047 = data_d1[111:104];
        6'd15: vec_data_047 = data_d1[119:112];
        6'd16: vec_data_047 = data_d1[127:120];
        6'd17: vec_data_047 = data_d1[135:128];
        6'd18: vec_data_047 = data_d1[143:136];
        6'd19: vec_data_047 = data_d1[151:144];
        6'd20: vec_data_047 = data_d1[159:152];
        6'd21: vec_data_047 = data_d1[167:160];
        6'd22: vec_data_047 = data_d1[175:168];
        6'd23: vec_data_047 = data_d1[183:176];
        6'd24: vec_data_047 = data_d1[191:184];
        6'd25: vec_data_047 = data_d1[199:192];
        6'd26: vec_data_047 = data_d1[207:200];
        6'd27: vec_data_047 = data_d1[215:208];
        6'd28: vec_data_047 = data_d1[223:216];
        6'd29: vec_data_047 = data_d1[231:224];
        6'd30: vec_data_047 = data_d1[239:232];
        6'd31: vec_data_047 = data_d1[247:240];
        6'd32: vec_data_047 = data_d1[255:248];
        6'd33: vec_data_047 = data_d1[263:256];
        6'd34: vec_data_047 = data_d1[271:264];
        6'd35: vec_data_047 = data_d1[279:272];
        6'd36: vec_data_047 = data_d1[287:280];
        6'd37: vec_data_047 = data_d1[295:288];
        6'd38: vec_data_047 = data_d1[303:296];
        6'd39: vec_data_047 = data_d1[311:304];
        6'd40: vec_data_047 = data_d1[319:312];
        6'd41: vec_data_047 = data_d1[327:320];
        6'd42: vec_data_047 = data_d1[335:328];
        6'd43: vec_data_047 = data_d1[343:336];
        6'd44: vec_data_047 = data_d1[351:344];
        6'd45: vec_data_047 = data_d1[359:352];
        6'd46: vec_data_047 = data_d1[367:360];
        6'd47: vec_data_047 = data_d1[375:368];
        6'd48: vec_data_047 = data_d1[383:376];
    endcase
end

always @(
  vec_sum_048_d1
  or data_d1
  ) begin
    vec_data_048 = 8'b0;
    case(vec_sum_048_d1)
        6'd1: vec_data_048 = data_d1[7:0];
        6'd2: vec_data_048 = data_d1[15:8];
        6'd3: vec_data_048 = data_d1[23:16];
        6'd4: vec_data_048 = data_d1[31:24];
        6'd5: vec_data_048 = data_d1[39:32];
        6'd6: vec_data_048 = data_d1[47:40];
        6'd7: vec_data_048 = data_d1[55:48];
        6'd8: vec_data_048 = data_d1[63:56];
        6'd9: vec_data_048 = data_d1[71:64];
        6'd10: vec_data_048 = data_d1[79:72];
        6'd11: vec_data_048 = data_d1[87:80];
        6'd12: vec_data_048 = data_d1[95:88];
        6'd13: vec_data_048 = data_d1[103:96];
        6'd14: vec_data_048 = data_d1[111:104];
        6'd15: vec_data_048 = data_d1[119:112];
        6'd16: vec_data_048 = data_d1[127:120];
        6'd17: vec_data_048 = data_d1[135:128];
        6'd18: vec_data_048 = data_d1[143:136];
        6'd19: vec_data_048 = data_d1[151:144];
        6'd20: vec_data_048 = data_d1[159:152];
        6'd21: vec_data_048 = data_d1[167:160];
        6'd22: vec_data_048 = data_d1[175:168];
        6'd23: vec_data_048 = data_d1[183:176];
        6'd24: vec_data_048 = data_d1[191:184];
        6'd25: vec_data_048 = data_d1[199:192];
        6'd26: vec_data_048 = data_d1[207:200];
        6'd27: vec_data_048 = data_d1[215:208];
        6'd28: vec_data_048 = data_d1[223:216];
        6'd29: vec_data_048 = data_d1[231:224];
        6'd30: vec_data_048 = data_d1[239:232];
        6'd31: vec_data_048 = data_d1[247:240];
        6'd32: vec_data_048 = data_d1[255:248];
        6'd33: vec_data_048 = data_d1[263:256];
        6'd34: vec_data_048 = data_d1[271:264];
        6'd35: vec_data_048 = data_d1[279:272];
        6'd36: vec_data_048 = data_d1[287:280];
        6'd37: vec_data_048 = data_d1[295:288];
        6'd38: vec_data_048 = data_d1[303:296];
        6'd39: vec_data_048 = data_d1[311:304];
        6'd40: vec_data_048 = data_d1[319:312];
        6'd41: vec_data_048 = data_d1[327:320];
        6'd42: vec_data_048 = data_d1[335:328];
        6'd43: vec_data_048 = data_d1[343:336];
        6'd44: vec_data_048 = data_d1[351:344];
        6'd45: vec_data_048 = data_d1[359:352];
        6'd46: vec_data_048 = data_d1[367:360];
        6'd47: vec_data_048 = data_d1[375:368];
        6'd48: vec_data_048 = data_d1[383:376];
        6'd49: vec_data_048 = data_d1[391:384];
    endcase
end

always @(
  vec_sum_049_d1
  or data_d1
  ) begin
    vec_data_049 = 8'b0;
    case(vec_sum_049_d1)
        6'd1: vec_data_049 = data_d1[7:0];
        6'd2: vec_data_049 = data_d1[15:8];
        6'd3: vec_data_049 = data_d1[23:16];
        6'd4: vec_data_049 = data_d1[31:24];
        6'd5: vec_data_049 = data_d1[39:32];
        6'd6: vec_data_049 = data_d1[47:40];
        6'd7: vec_data_049 = data_d1[55:48];
        6'd8: vec_data_049 = data_d1[63:56];
        6'd9: vec_data_049 = data_d1[71:64];
        6'd10: vec_data_049 = data_d1[79:72];
        6'd11: vec_data_049 = data_d1[87:80];
        6'd12: vec_data_049 = data_d1[95:88];
        6'd13: vec_data_049 = data_d1[103:96];
        6'd14: vec_data_049 = data_d1[111:104];
        6'd15: vec_data_049 = data_d1[119:112];
        6'd16: vec_data_049 = data_d1[127:120];
        6'd17: vec_data_049 = data_d1[135:128];
        6'd18: vec_data_049 = data_d1[143:136];
        6'd19: vec_data_049 = data_d1[151:144];
        6'd20: vec_data_049 = data_d1[159:152];
        6'd21: vec_data_049 = data_d1[167:160];
        6'd22: vec_data_049 = data_d1[175:168];
        6'd23: vec_data_049 = data_d1[183:176];
        6'd24: vec_data_049 = data_d1[191:184];
        6'd25: vec_data_049 = data_d1[199:192];
        6'd26: vec_data_049 = data_d1[207:200];
        6'd27: vec_data_049 = data_d1[215:208];
        6'd28: vec_data_049 = data_d1[223:216];
        6'd29: vec_data_049 = data_d1[231:224];
        6'd30: vec_data_049 = data_d1[239:232];
        6'd31: vec_data_049 = data_d1[247:240];
        6'd32: vec_data_049 = data_d1[255:248];
        6'd33: vec_data_049 = data_d1[263:256];
        6'd34: vec_data_049 = data_d1[271:264];
        6'd35: vec_data_049 = data_d1[279:272];
        6'd36: vec_data_049 = data_d1[287:280];
        6'd37: vec_data_049 = data_d1[295:288];
        6'd38: vec_data_049 = data_d1[303:296];
        6'd39: vec_data_049 = data_d1[311:304];
        6'd40: vec_data_049 = data_d1[319:312];
        6'd41: vec_data_049 = data_d1[327:320];
        6'd42: vec_data_049 = data_d1[335:328];
        6'd43: vec_data_049 = data_d1[343:336];
        6'd44: vec_data_049 = data_d1[351:344];
        6'd45: vec_data_049 = data_d1[359:352];
        6'd46: vec_data_049 = data_d1[367:360];
        6'd47: vec_data_049 = data_d1[375:368];
        6'd48: vec_data_049 = data_d1[383:376];
        6'd49: vec_data_049 = data_d1[391:384];
        6'd50: vec_data_049 = data_d1[399:392];
    endcase
end

always @(
  vec_sum_050_d1
  or data_d1
  ) begin
    vec_data_050 = 8'b0;
    case(vec_sum_050_d1)
        6'd1: vec_data_050 = data_d1[7:0];
        6'd2: vec_data_050 = data_d1[15:8];
        6'd3: vec_data_050 = data_d1[23:16];
        6'd4: vec_data_050 = data_d1[31:24];
        6'd5: vec_data_050 = data_d1[39:32];
        6'd6: vec_data_050 = data_d1[47:40];
        6'd7: vec_data_050 = data_d1[55:48];
        6'd8: vec_data_050 = data_d1[63:56];
        6'd9: vec_data_050 = data_d1[71:64];
        6'd10: vec_data_050 = data_d1[79:72];
        6'd11: vec_data_050 = data_d1[87:80];
        6'd12: vec_data_050 = data_d1[95:88];
        6'd13: vec_data_050 = data_d1[103:96];
        6'd14: vec_data_050 = data_d1[111:104];
        6'd15: vec_data_050 = data_d1[119:112];
        6'd16: vec_data_050 = data_d1[127:120];
        6'd17: vec_data_050 = data_d1[135:128];
        6'd18: vec_data_050 = data_d1[143:136];
        6'd19: vec_data_050 = data_d1[151:144];
        6'd20: vec_data_050 = data_d1[159:152];
        6'd21: vec_data_050 = data_d1[167:160];
        6'd22: vec_data_050 = data_d1[175:168];
        6'd23: vec_data_050 = data_d1[183:176];
        6'd24: vec_data_050 = data_d1[191:184];
        6'd25: vec_data_050 = data_d1[199:192];
        6'd26: vec_data_050 = data_d1[207:200];
        6'd27: vec_data_050 = data_d1[215:208];
        6'd28: vec_data_050 = data_d1[223:216];
        6'd29: vec_data_050 = data_d1[231:224];
        6'd30: vec_data_050 = data_d1[239:232];
        6'd31: vec_data_050 = data_d1[247:240];
        6'd32: vec_data_050 = data_d1[255:248];
        6'd33: vec_data_050 = data_d1[263:256];
        6'd34: vec_data_050 = data_d1[271:264];
        6'd35: vec_data_050 = data_d1[279:272];
        6'd36: vec_data_050 = data_d1[287:280];
        6'd37: vec_data_050 = data_d1[295:288];
        6'd38: vec_data_050 = data_d1[303:296];
        6'd39: vec_data_050 = data_d1[311:304];
        6'd40: vec_data_050 = data_d1[319:312];
        6'd41: vec_data_050 = data_d1[327:320];
        6'd42: vec_data_050 = data_d1[335:328];
        6'd43: vec_data_050 = data_d1[343:336];
        6'd44: vec_data_050 = data_d1[351:344];
        6'd45: vec_data_050 = data_d1[359:352];
        6'd46: vec_data_050 = data_d1[367:360];
        6'd47: vec_data_050 = data_d1[375:368];
        6'd48: vec_data_050 = data_d1[383:376];
        6'd49: vec_data_050 = data_d1[391:384];
        6'd50: vec_data_050 = data_d1[399:392];
        6'd51: vec_data_050 = data_d1[407:400];
    endcase
end

always @(
  vec_sum_051_d1
  or data_d1
  ) begin
    vec_data_051 = 8'b0;
    case(vec_sum_051_d1)
        6'd1: vec_data_051 = data_d1[7:0];
        6'd2: vec_data_051 = data_d1[15:8];
        6'd3: vec_data_051 = data_d1[23:16];
        6'd4: vec_data_051 = data_d1[31:24];
        6'd5: vec_data_051 = data_d1[39:32];
        6'd6: vec_data_051 = data_d1[47:40];
        6'd7: vec_data_051 = data_d1[55:48];
        6'd8: vec_data_051 = data_d1[63:56];
        6'd9: vec_data_051 = data_d1[71:64];
        6'd10: vec_data_051 = data_d1[79:72];
        6'd11: vec_data_051 = data_d1[87:80];
        6'd12: vec_data_051 = data_d1[95:88];
        6'd13: vec_data_051 = data_d1[103:96];
        6'd14: vec_data_051 = data_d1[111:104];
        6'd15: vec_data_051 = data_d1[119:112];
        6'd16: vec_data_051 = data_d1[127:120];
        6'd17: vec_data_051 = data_d1[135:128];
        6'd18: vec_data_051 = data_d1[143:136];
        6'd19: vec_data_051 = data_d1[151:144];
        6'd20: vec_data_051 = data_d1[159:152];
        6'd21: vec_data_051 = data_d1[167:160];
        6'd22: vec_data_051 = data_d1[175:168];
        6'd23: vec_data_051 = data_d1[183:176];
        6'd24: vec_data_051 = data_d1[191:184];
        6'd25: vec_data_051 = data_d1[199:192];
        6'd26: vec_data_051 = data_d1[207:200];
        6'd27: vec_data_051 = data_d1[215:208];
        6'd28: vec_data_051 = data_d1[223:216];
        6'd29: vec_data_051 = data_d1[231:224];
        6'd30: vec_data_051 = data_d1[239:232];
        6'd31: vec_data_051 = data_d1[247:240];
        6'd32: vec_data_051 = data_d1[255:248];
        6'd33: vec_data_051 = data_d1[263:256];
        6'd34: vec_data_051 = data_d1[271:264];
        6'd35: vec_data_051 = data_d1[279:272];
        6'd36: vec_data_051 = data_d1[287:280];
        6'd37: vec_data_051 = data_d1[295:288];
        6'd38: vec_data_051 = data_d1[303:296];
        6'd39: vec_data_051 = data_d1[311:304];
        6'd40: vec_data_051 = data_d1[319:312];
        6'd41: vec_data_051 = data_d1[327:320];
        6'd42: vec_data_051 = data_d1[335:328];
        6'd43: vec_data_051 = data_d1[343:336];
        6'd44: vec_data_051 = data_d1[351:344];
        6'd45: vec_data_051 = data_d1[359:352];
        6'd46: vec_data_051 = data_d1[367:360];
        6'd47: vec_data_051 = data_d1[375:368];
        6'd48: vec_data_051 = data_d1[383:376];
        6'd49: vec_data_051 = data_d1[391:384];
        6'd50: vec_data_051 = data_d1[399:392];
        6'd51: vec_data_051 = data_d1[407:400];
        6'd52: vec_data_051 = data_d1[415:408];
    endcase
end

always @(
  vec_sum_052_d1
  or data_d1
  ) begin
    vec_data_052 = 8'b0;
    case(vec_sum_052_d1)
        6'd1: vec_data_052 = data_d1[7:0];
        6'd2: vec_data_052 = data_d1[15:8];
        6'd3: vec_data_052 = data_d1[23:16];
        6'd4: vec_data_052 = data_d1[31:24];
        6'd5: vec_data_052 = data_d1[39:32];
        6'd6: vec_data_052 = data_d1[47:40];
        6'd7: vec_data_052 = data_d1[55:48];
        6'd8: vec_data_052 = data_d1[63:56];
        6'd9: vec_data_052 = data_d1[71:64];
        6'd10: vec_data_052 = data_d1[79:72];
        6'd11: vec_data_052 = data_d1[87:80];
        6'd12: vec_data_052 = data_d1[95:88];
        6'd13: vec_data_052 = data_d1[103:96];
        6'd14: vec_data_052 = data_d1[111:104];
        6'd15: vec_data_052 = data_d1[119:112];
        6'd16: vec_data_052 = data_d1[127:120];
        6'd17: vec_data_052 = data_d1[135:128];
        6'd18: vec_data_052 = data_d1[143:136];
        6'd19: vec_data_052 = data_d1[151:144];
        6'd20: vec_data_052 = data_d1[159:152];
        6'd21: vec_data_052 = data_d1[167:160];
        6'd22: vec_data_052 = data_d1[175:168];
        6'd23: vec_data_052 = data_d1[183:176];
        6'd24: vec_data_052 = data_d1[191:184];
        6'd25: vec_data_052 = data_d1[199:192];
        6'd26: vec_data_052 = data_d1[207:200];
        6'd27: vec_data_052 = data_d1[215:208];
        6'd28: vec_data_052 = data_d1[223:216];
        6'd29: vec_data_052 = data_d1[231:224];
        6'd30: vec_data_052 = data_d1[239:232];
        6'd31: vec_data_052 = data_d1[247:240];
        6'd32: vec_data_052 = data_d1[255:248];
        6'd33: vec_data_052 = data_d1[263:256];
        6'd34: vec_data_052 = data_d1[271:264];
        6'd35: vec_data_052 = data_d1[279:272];
        6'd36: vec_data_052 = data_d1[287:280];
        6'd37: vec_data_052 = data_d1[295:288];
        6'd38: vec_data_052 = data_d1[303:296];
        6'd39: vec_data_052 = data_d1[311:304];
        6'd40: vec_data_052 = data_d1[319:312];
        6'd41: vec_data_052 = data_d1[327:320];
        6'd42: vec_data_052 = data_d1[335:328];
        6'd43: vec_data_052 = data_d1[343:336];
        6'd44: vec_data_052 = data_d1[351:344];
        6'd45: vec_data_052 = data_d1[359:352];
        6'd46: vec_data_052 = data_d1[367:360];
        6'd47: vec_data_052 = data_d1[375:368];
        6'd48: vec_data_052 = data_d1[383:376];
        6'd49: vec_data_052 = data_d1[391:384];
        6'd50: vec_data_052 = data_d1[399:392];
        6'd51: vec_data_052 = data_d1[407:400];
        6'd52: vec_data_052 = data_d1[415:408];
        6'd53: vec_data_052 = data_d1[423:416];
    endcase
end

always @(
  vec_sum_053_d1
  or data_d1
  ) begin
    vec_data_053 = 8'b0;
    case(vec_sum_053_d1)
        6'd1: vec_data_053 = data_d1[7:0];
        6'd2: vec_data_053 = data_d1[15:8];
        6'd3: vec_data_053 = data_d1[23:16];
        6'd4: vec_data_053 = data_d1[31:24];
        6'd5: vec_data_053 = data_d1[39:32];
        6'd6: vec_data_053 = data_d1[47:40];
        6'd7: vec_data_053 = data_d1[55:48];
        6'd8: vec_data_053 = data_d1[63:56];
        6'd9: vec_data_053 = data_d1[71:64];
        6'd10: vec_data_053 = data_d1[79:72];
        6'd11: vec_data_053 = data_d1[87:80];
        6'd12: vec_data_053 = data_d1[95:88];
        6'd13: vec_data_053 = data_d1[103:96];
        6'd14: vec_data_053 = data_d1[111:104];
        6'd15: vec_data_053 = data_d1[119:112];
        6'd16: vec_data_053 = data_d1[127:120];
        6'd17: vec_data_053 = data_d1[135:128];
        6'd18: vec_data_053 = data_d1[143:136];
        6'd19: vec_data_053 = data_d1[151:144];
        6'd20: vec_data_053 = data_d1[159:152];
        6'd21: vec_data_053 = data_d1[167:160];
        6'd22: vec_data_053 = data_d1[175:168];
        6'd23: vec_data_053 = data_d1[183:176];
        6'd24: vec_data_053 = data_d1[191:184];
        6'd25: vec_data_053 = data_d1[199:192];
        6'd26: vec_data_053 = data_d1[207:200];
        6'd27: vec_data_053 = data_d1[215:208];
        6'd28: vec_data_053 = data_d1[223:216];
        6'd29: vec_data_053 = data_d1[231:224];
        6'd30: vec_data_053 = data_d1[239:232];
        6'd31: vec_data_053 = data_d1[247:240];
        6'd32: vec_data_053 = data_d1[255:248];
        6'd33: vec_data_053 = data_d1[263:256];
        6'd34: vec_data_053 = data_d1[271:264];
        6'd35: vec_data_053 = data_d1[279:272];
        6'd36: vec_data_053 = data_d1[287:280];
        6'd37: vec_data_053 = data_d1[295:288];
        6'd38: vec_data_053 = data_d1[303:296];
        6'd39: vec_data_053 = data_d1[311:304];
        6'd40: vec_data_053 = data_d1[319:312];
        6'd41: vec_data_053 = data_d1[327:320];
        6'd42: vec_data_053 = data_d1[335:328];
        6'd43: vec_data_053 = data_d1[343:336];
        6'd44: vec_data_053 = data_d1[351:344];
        6'd45: vec_data_053 = data_d1[359:352];
        6'd46: vec_data_053 = data_d1[367:360];
        6'd47: vec_data_053 = data_d1[375:368];
        6'd48: vec_data_053 = data_d1[383:376];
        6'd49: vec_data_053 = data_d1[391:384];
        6'd50: vec_data_053 = data_d1[399:392];
        6'd51: vec_data_053 = data_d1[407:400];
        6'd52: vec_data_053 = data_d1[415:408];
        6'd53: vec_data_053 = data_d1[423:416];
        6'd54: vec_data_053 = data_d1[431:424];
    endcase
end

always @(
  vec_sum_054_d1
  or data_d1
  ) begin
    vec_data_054 = 8'b0;
    case(vec_sum_054_d1)
        6'd1: vec_data_054 = data_d1[7:0];
        6'd2: vec_data_054 = data_d1[15:8];
        6'd3: vec_data_054 = data_d1[23:16];
        6'd4: vec_data_054 = data_d1[31:24];
        6'd5: vec_data_054 = data_d1[39:32];
        6'd6: vec_data_054 = data_d1[47:40];
        6'd7: vec_data_054 = data_d1[55:48];
        6'd8: vec_data_054 = data_d1[63:56];
        6'd9: vec_data_054 = data_d1[71:64];
        6'd10: vec_data_054 = data_d1[79:72];
        6'd11: vec_data_054 = data_d1[87:80];
        6'd12: vec_data_054 = data_d1[95:88];
        6'd13: vec_data_054 = data_d1[103:96];
        6'd14: vec_data_054 = data_d1[111:104];
        6'd15: vec_data_054 = data_d1[119:112];
        6'd16: vec_data_054 = data_d1[127:120];
        6'd17: vec_data_054 = data_d1[135:128];
        6'd18: vec_data_054 = data_d1[143:136];
        6'd19: vec_data_054 = data_d1[151:144];
        6'd20: vec_data_054 = data_d1[159:152];
        6'd21: vec_data_054 = data_d1[167:160];
        6'd22: vec_data_054 = data_d1[175:168];
        6'd23: vec_data_054 = data_d1[183:176];
        6'd24: vec_data_054 = data_d1[191:184];
        6'd25: vec_data_054 = data_d1[199:192];
        6'd26: vec_data_054 = data_d1[207:200];
        6'd27: vec_data_054 = data_d1[215:208];
        6'd28: vec_data_054 = data_d1[223:216];
        6'd29: vec_data_054 = data_d1[231:224];
        6'd30: vec_data_054 = data_d1[239:232];
        6'd31: vec_data_054 = data_d1[247:240];
        6'd32: vec_data_054 = data_d1[255:248];
        6'd33: vec_data_054 = data_d1[263:256];
        6'd34: vec_data_054 = data_d1[271:264];
        6'd35: vec_data_054 = data_d1[279:272];
        6'd36: vec_data_054 = data_d1[287:280];
        6'd37: vec_data_054 = data_d1[295:288];
        6'd38: vec_data_054 = data_d1[303:296];
        6'd39: vec_data_054 = data_d1[311:304];
        6'd40: vec_data_054 = data_d1[319:312];
        6'd41: vec_data_054 = data_d1[327:320];
        6'd42: vec_data_054 = data_d1[335:328];
        6'd43: vec_data_054 = data_d1[343:336];
        6'd44: vec_data_054 = data_d1[351:344];
        6'd45: vec_data_054 = data_d1[359:352];
        6'd46: vec_data_054 = data_d1[367:360];
        6'd47: vec_data_054 = data_d1[375:368];
        6'd48: vec_data_054 = data_d1[383:376];
        6'd49: vec_data_054 = data_d1[391:384];
        6'd50: vec_data_054 = data_d1[399:392];
        6'd51: vec_data_054 = data_d1[407:400];
        6'd52: vec_data_054 = data_d1[415:408];
        6'd53: vec_data_054 = data_d1[423:416];
        6'd54: vec_data_054 = data_d1[431:424];
        6'd55: vec_data_054 = data_d1[439:432];
    endcase
end

always @(
  vec_sum_055_d1
  or data_d1
  ) begin
    vec_data_055 = 8'b0;
    case(vec_sum_055_d1)
        6'd1: vec_data_055 = data_d1[7:0];
        6'd2: vec_data_055 = data_d1[15:8];
        6'd3: vec_data_055 = data_d1[23:16];
        6'd4: vec_data_055 = data_d1[31:24];
        6'd5: vec_data_055 = data_d1[39:32];
        6'd6: vec_data_055 = data_d1[47:40];
        6'd7: vec_data_055 = data_d1[55:48];
        6'd8: vec_data_055 = data_d1[63:56];
        6'd9: vec_data_055 = data_d1[71:64];
        6'd10: vec_data_055 = data_d1[79:72];
        6'd11: vec_data_055 = data_d1[87:80];
        6'd12: vec_data_055 = data_d1[95:88];
        6'd13: vec_data_055 = data_d1[103:96];
        6'd14: vec_data_055 = data_d1[111:104];
        6'd15: vec_data_055 = data_d1[119:112];
        6'd16: vec_data_055 = data_d1[127:120];
        6'd17: vec_data_055 = data_d1[135:128];
        6'd18: vec_data_055 = data_d1[143:136];
        6'd19: vec_data_055 = data_d1[151:144];
        6'd20: vec_data_055 = data_d1[159:152];
        6'd21: vec_data_055 = data_d1[167:160];
        6'd22: vec_data_055 = data_d1[175:168];
        6'd23: vec_data_055 = data_d1[183:176];
        6'd24: vec_data_055 = data_d1[191:184];
        6'd25: vec_data_055 = data_d1[199:192];
        6'd26: vec_data_055 = data_d1[207:200];
        6'd27: vec_data_055 = data_d1[215:208];
        6'd28: vec_data_055 = data_d1[223:216];
        6'd29: vec_data_055 = data_d1[231:224];
        6'd30: vec_data_055 = data_d1[239:232];
        6'd31: vec_data_055 = data_d1[247:240];
        6'd32: vec_data_055 = data_d1[255:248];
        6'd33: vec_data_055 = data_d1[263:256];
        6'd34: vec_data_055 = data_d1[271:264];
        6'd35: vec_data_055 = data_d1[279:272];
        6'd36: vec_data_055 = data_d1[287:280];
        6'd37: vec_data_055 = data_d1[295:288];
        6'd38: vec_data_055 = data_d1[303:296];
        6'd39: vec_data_055 = data_d1[311:304];
        6'd40: vec_data_055 = data_d1[319:312];
        6'd41: vec_data_055 = data_d1[327:320];
        6'd42: vec_data_055 = data_d1[335:328];
        6'd43: vec_data_055 = data_d1[343:336];
        6'd44: vec_data_055 = data_d1[351:344];
        6'd45: vec_data_055 = data_d1[359:352];
        6'd46: vec_data_055 = data_d1[367:360];
        6'd47: vec_data_055 = data_d1[375:368];
        6'd48: vec_data_055 = data_d1[383:376];
        6'd49: vec_data_055 = data_d1[391:384];
        6'd50: vec_data_055 = data_d1[399:392];
        6'd51: vec_data_055 = data_d1[407:400];
        6'd52: vec_data_055 = data_d1[415:408];
        6'd53: vec_data_055 = data_d1[423:416];
        6'd54: vec_data_055 = data_d1[431:424];
        6'd55: vec_data_055 = data_d1[439:432];
        6'd56: vec_data_055 = data_d1[447:440];
    endcase
end

always @(
  vec_sum_056_d1
  or data_d1
  ) begin
    vec_data_056 = 8'b0;
    case(vec_sum_056_d1)
        6'd1: vec_data_056 = data_d1[7:0];
        6'd2: vec_data_056 = data_d1[15:8];
        6'd3: vec_data_056 = data_d1[23:16];
        6'd4: vec_data_056 = data_d1[31:24];
        6'd5: vec_data_056 = data_d1[39:32];
        6'd6: vec_data_056 = data_d1[47:40];
        6'd7: vec_data_056 = data_d1[55:48];
        6'd8: vec_data_056 = data_d1[63:56];
        6'd9: vec_data_056 = data_d1[71:64];
        6'd10: vec_data_056 = data_d1[79:72];
        6'd11: vec_data_056 = data_d1[87:80];
        6'd12: vec_data_056 = data_d1[95:88];
        6'd13: vec_data_056 = data_d1[103:96];
        6'd14: vec_data_056 = data_d1[111:104];
        6'd15: vec_data_056 = data_d1[119:112];
        6'd16: vec_data_056 = data_d1[127:120];
        6'd17: vec_data_056 = data_d1[135:128];
        6'd18: vec_data_056 = data_d1[143:136];
        6'd19: vec_data_056 = data_d1[151:144];
        6'd20: vec_data_056 = data_d1[159:152];
        6'd21: vec_data_056 = data_d1[167:160];
        6'd22: vec_data_056 = data_d1[175:168];
        6'd23: vec_data_056 = data_d1[183:176];
        6'd24: vec_data_056 = data_d1[191:184];
        6'd25: vec_data_056 = data_d1[199:192];
        6'd26: vec_data_056 = data_d1[207:200];
        6'd27: vec_data_056 = data_d1[215:208];
        6'd28: vec_data_056 = data_d1[223:216];
        6'd29: vec_data_056 = data_d1[231:224];
        6'd30: vec_data_056 = data_d1[239:232];
        6'd31: vec_data_056 = data_d1[247:240];
        6'd32: vec_data_056 = data_d1[255:248];
        6'd33: vec_data_056 = data_d1[263:256];
        6'd34: vec_data_056 = data_d1[271:264];
        6'd35: vec_data_056 = data_d1[279:272];
        6'd36: vec_data_056 = data_d1[287:280];
        6'd37: vec_data_056 = data_d1[295:288];
        6'd38: vec_data_056 = data_d1[303:296];
        6'd39: vec_data_056 = data_d1[311:304];
        6'd40: vec_data_056 = data_d1[319:312];
        6'd41: vec_data_056 = data_d1[327:320];
        6'd42: vec_data_056 = data_d1[335:328];
        6'd43: vec_data_056 = data_d1[343:336];
        6'd44: vec_data_056 = data_d1[351:344];
        6'd45: vec_data_056 = data_d1[359:352];
        6'd46: vec_data_056 = data_d1[367:360];
        6'd47: vec_data_056 = data_d1[375:368];
        6'd48: vec_data_056 = data_d1[383:376];
        6'd49: vec_data_056 = data_d1[391:384];
        6'd50: vec_data_056 = data_d1[399:392];
        6'd51: vec_data_056 = data_d1[407:400];
        6'd52: vec_data_056 = data_d1[415:408];
        6'd53: vec_data_056 = data_d1[423:416];
        6'd54: vec_data_056 = data_d1[431:424];
        6'd55: vec_data_056 = data_d1[439:432];
        6'd56: vec_data_056 = data_d1[447:440];
        6'd57: vec_data_056 = data_d1[455:448];
    endcase
end

always @(
  vec_sum_057_d1
  or data_d1
  ) begin
    vec_data_057 = 8'b0;
    case(vec_sum_057_d1)
        6'd1: vec_data_057 = data_d1[7:0];
        6'd2: vec_data_057 = data_d1[15:8];
        6'd3: vec_data_057 = data_d1[23:16];
        6'd4: vec_data_057 = data_d1[31:24];
        6'd5: vec_data_057 = data_d1[39:32];
        6'd6: vec_data_057 = data_d1[47:40];
        6'd7: vec_data_057 = data_d1[55:48];
        6'd8: vec_data_057 = data_d1[63:56];
        6'd9: vec_data_057 = data_d1[71:64];
        6'd10: vec_data_057 = data_d1[79:72];
        6'd11: vec_data_057 = data_d1[87:80];
        6'd12: vec_data_057 = data_d1[95:88];
        6'd13: vec_data_057 = data_d1[103:96];
        6'd14: vec_data_057 = data_d1[111:104];
        6'd15: vec_data_057 = data_d1[119:112];
        6'd16: vec_data_057 = data_d1[127:120];
        6'd17: vec_data_057 = data_d1[135:128];
        6'd18: vec_data_057 = data_d1[143:136];
        6'd19: vec_data_057 = data_d1[151:144];
        6'd20: vec_data_057 = data_d1[159:152];
        6'd21: vec_data_057 = data_d1[167:160];
        6'd22: vec_data_057 = data_d1[175:168];
        6'd23: vec_data_057 = data_d1[183:176];
        6'd24: vec_data_057 = data_d1[191:184];
        6'd25: vec_data_057 = data_d1[199:192];
        6'd26: vec_data_057 = data_d1[207:200];
        6'd27: vec_data_057 = data_d1[215:208];
        6'd28: vec_data_057 = data_d1[223:216];
        6'd29: vec_data_057 = data_d1[231:224];
        6'd30: vec_data_057 = data_d1[239:232];
        6'd31: vec_data_057 = data_d1[247:240];
        6'd32: vec_data_057 = data_d1[255:248];
        6'd33: vec_data_057 = data_d1[263:256];
        6'd34: vec_data_057 = data_d1[271:264];
        6'd35: vec_data_057 = data_d1[279:272];
        6'd36: vec_data_057 = data_d1[287:280];
        6'd37: vec_data_057 = data_d1[295:288];
        6'd38: vec_data_057 = data_d1[303:296];
        6'd39: vec_data_057 = data_d1[311:304];
        6'd40: vec_data_057 = data_d1[319:312];
        6'd41: vec_data_057 = data_d1[327:320];
        6'd42: vec_data_057 = data_d1[335:328];
        6'd43: vec_data_057 = data_d1[343:336];
        6'd44: vec_data_057 = data_d1[351:344];
        6'd45: vec_data_057 = data_d1[359:352];
        6'd46: vec_data_057 = data_d1[367:360];
        6'd47: vec_data_057 = data_d1[375:368];
        6'd48: vec_data_057 = data_d1[383:376];
        6'd49: vec_data_057 = data_d1[391:384];
        6'd50: vec_data_057 = data_d1[399:392];
        6'd51: vec_data_057 = data_d1[407:400];
        6'd52: vec_data_057 = data_d1[415:408];
        6'd53: vec_data_057 = data_d1[423:416];
        6'd54: vec_data_057 = data_d1[431:424];
        6'd55: vec_data_057 = data_d1[439:432];
        6'd56: vec_data_057 = data_d1[447:440];
        6'd57: vec_data_057 = data_d1[455:448];
        6'd58: vec_data_057 = data_d1[463:456];
    endcase
end

always @(
  vec_sum_058_d1
  or data_d1
  ) begin
    vec_data_058 = 8'b0;
    case(vec_sum_058_d1)
        6'd1: vec_data_058 = data_d1[7:0];
        6'd2: vec_data_058 = data_d1[15:8];
        6'd3: vec_data_058 = data_d1[23:16];
        6'd4: vec_data_058 = data_d1[31:24];
        6'd5: vec_data_058 = data_d1[39:32];
        6'd6: vec_data_058 = data_d1[47:40];
        6'd7: vec_data_058 = data_d1[55:48];
        6'd8: vec_data_058 = data_d1[63:56];
        6'd9: vec_data_058 = data_d1[71:64];
        6'd10: vec_data_058 = data_d1[79:72];
        6'd11: vec_data_058 = data_d1[87:80];
        6'd12: vec_data_058 = data_d1[95:88];
        6'd13: vec_data_058 = data_d1[103:96];
        6'd14: vec_data_058 = data_d1[111:104];
        6'd15: vec_data_058 = data_d1[119:112];
        6'd16: vec_data_058 = data_d1[127:120];
        6'd17: vec_data_058 = data_d1[135:128];
        6'd18: vec_data_058 = data_d1[143:136];
        6'd19: vec_data_058 = data_d1[151:144];
        6'd20: vec_data_058 = data_d1[159:152];
        6'd21: vec_data_058 = data_d1[167:160];
        6'd22: vec_data_058 = data_d1[175:168];
        6'd23: vec_data_058 = data_d1[183:176];
        6'd24: vec_data_058 = data_d1[191:184];
        6'd25: vec_data_058 = data_d1[199:192];
        6'd26: vec_data_058 = data_d1[207:200];
        6'd27: vec_data_058 = data_d1[215:208];
        6'd28: vec_data_058 = data_d1[223:216];
        6'd29: vec_data_058 = data_d1[231:224];
        6'd30: vec_data_058 = data_d1[239:232];
        6'd31: vec_data_058 = data_d1[247:240];
        6'd32: vec_data_058 = data_d1[255:248];
        6'd33: vec_data_058 = data_d1[263:256];
        6'd34: vec_data_058 = data_d1[271:264];
        6'd35: vec_data_058 = data_d1[279:272];
        6'd36: vec_data_058 = data_d1[287:280];
        6'd37: vec_data_058 = data_d1[295:288];
        6'd38: vec_data_058 = data_d1[303:296];
        6'd39: vec_data_058 = data_d1[311:304];
        6'd40: vec_data_058 = data_d1[319:312];
        6'd41: vec_data_058 = data_d1[327:320];
        6'd42: vec_data_058 = data_d1[335:328];
        6'd43: vec_data_058 = data_d1[343:336];
        6'd44: vec_data_058 = data_d1[351:344];
        6'd45: vec_data_058 = data_d1[359:352];
        6'd46: vec_data_058 = data_d1[367:360];
        6'd47: vec_data_058 = data_d1[375:368];
        6'd48: vec_data_058 = data_d1[383:376];
        6'd49: vec_data_058 = data_d1[391:384];
        6'd50: vec_data_058 = data_d1[399:392];
        6'd51: vec_data_058 = data_d1[407:400];
        6'd52: vec_data_058 = data_d1[415:408];
        6'd53: vec_data_058 = data_d1[423:416];
        6'd54: vec_data_058 = data_d1[431:424];
        6'd55: vec_data_058 = data_d1[439:432];
        6'd56: vec_data_058 = data_d1[447:440];
        6'd57: vec_data_058 = data_d1[455:448];
        6'd58: vec_data_058 = data_d1[463:456];
        6'd59: vec_data_058 = data_d1[471:464];
    endcase
end

always @(
  vec_sum_059_d1
  or data_d1
  ) begin
    vec_data_059 = 8'b0;
    case(vec_sum_059_d1)
        6'd1: vec_data_059 = data_d1[7:0];
        6'd2: vec_data_059 = data_d1[15:8];
        6'd3: vec_data_059 = data_d1[23:16];
        6'd4: vec_data_059 = data_d1[31:24];
        6'd5: vec_data_059 = data_d1[39:32];
        6'd6: vec_data_059 = data_d1[47:40];
        6'd7: vec_data_059 = data_d1[55:48];
        6'd8: vec_data_059 = data_d1[63:56];
        6'd9: vec_data_059 = data_d1[71:64];
        6'd10: vec_data_059 = data_d1[79:72];
        6'd11: vec_data_059 = data_d1[87:80];
        6'd12: vec_data_059 = data_d1[95:88];
        6'd13: vec_data_059 = data_d1[103:96];
        6'd14: vec_data_059 = data_d1[111:104];
        6'd15: vec_data_059 = data_d1[119:112];
        6'd16: vec_data_059 = data_d1[127:120];
        6'd17: vec_data_059 = data_d1[135:128];
        6'd18: vec_data_059 = data_d1[143:136];
        6'd19: vec_data_059 = data_d1[151:144];
        6'd20: vec_data_059 = data_d1[159:152];
        6'd21: vec_data_059 = data_d1[167:160];
        6'd22: vec_data_059 = data_d1[175:168];
        6'd23: vec_data_059 = data_d1[183:176];
        6'd24: vec_data_059 = data_d1[191:184];
        6'd25: vec_data_059 = data_d1[199:192];
        6'd26: vec_data_059 = data_d1[207:200];
        6'd27: vec_data_059 = data_d1[215:208];
        6'd28: vec_data_059 = data_d1[223:216];
        6'd29: vec_data_059 = data_d1[231:224];
        6'd30: vec_data_059 = data_d1[239:232];
        6'd31: vec_data_059 = data_d1[247:240];
        6'd32: vec_data_059 = data_d1[255:248];
        6'd33: vec_data_059 = data_d1[263:256];
        6'd34: vec_data_059 = data_d1[271:264];
        6'd35: vec_data_059 = data_d1[279:272];
        6'd36: vec_data_059 = data_d1[287:280];
        6'd37: vec_data_059 = data_d1[295:288];
        6'd38: vec_data_059 = data_d1[303:296];
        6'd39: vec_data_059 = data_d1[311:304];
        6'd40: vec_data_059 = data_d1[319:312];
        6'd41: vec_data_059 = data_d1[327:320];
        6'd42: vec_data_059 = data_d1[335:328];
        6'd43: vec_data_059 = data_d1[343:336];
        6'd44: vec_data_059 = data_d1[351:344];
        6'd45: vec_data_059 = data_d1[359:352];
        6'd46: vec_data_059 = data_d1[367:360];
        6'd47: vec_data_059 = data_d1[375:368];
        6'd48: vec_data_059 = data_d1[383:376];
        6'd49: vec_data_059 = data_d1[391:384];
        6'd50: vec_data_059 = data_d1[399:392];
        6'd51: vec_data_059 = data_d1[407:400];
        6'd52: vec_data_059 = data_d1[415:408];
        6'd53: vec_data_059 = data_d1[423:416];
        6'd54: vec_data_059 = data_d1[431:424];
        6'd55: vec_data_059 = data_d1[439:432];
        6'd56: vec_data_059 = data_d1[447:440];
        6'd57: vec_data_059 = data_d1[455:448];
        6'd58: vec_data_059 = data_d1[463:456];
        6'd59: vec_data_059 = data_d1[471:464];
        6'd60: vec_data_059 = data_d1[479:472];
    endcase
end

always @(
  vec_sum_060_d1
  or data_d1
  ) begin
    vec_data_060 = 8'b0;
    case(vec_sum_060_d1)
        6'd1: vec_data_060 = data_d1[7:0];
        6'd2: vec_data_060 = data_d1[15:8];
        6'd3: vec_data_060 = data_d1[23:16];
        6'd4: vec_data_060 = data_d1[31:24];
        6'd5: vec_data_060 = data_d1[39:32];
        6'd6: vec_data_060 = data_d1[47:40];
        6'd7: vec_data_060 = data_d1[55:48];
        6'd8: vec_data_060 = data_d1[63:56];
        6'd9: vec_data_060 = data_d1[71:64];
        6'd10: vec_data_060 = data_d1[79:72];
        6'd11: vec_data_060 = data_d1[87:80];
        6'd12: vec_data_060 = data_d1[95:88];
        6'd13: vec_data_060 = data_d1[103:96];
        6'd14: vec_data_060 = data_d1[111:104];
        6'd15: vec_data_060 = data_d1[119:112];
        6'd16: vec_data_060 = data_d1[127:120];
        6'd17: vec_data_060 = data_d1[135:128];
        6'd18: vec_data_060 = data_d1[143:136];
        6'd19: vec_data_060 = data_d1[151:144];
        6'd20: vec_data_060 = data_d1[159:152];
        6'd21: vec_data_060 = data_d1[167:160];
        6'd22: vec_data_060 = data_d1[175:168];
        6'd23: vec_data_060 = data_d1[183:176];
        6'd24: vec_data_060 = data_d1[191:184];
        6'd25: vec_data_060 = data_d1[199:192];
        6'd26: vec_data_060 = data_d1[207:200];
        6'd27: vec_data_060 = data_d1[215:208];
        6'd28: vec_data_060 = data_d1[223:216];
        6'd29: vec_data_060 = data_d1[231:224];
        6'd30: vec_data_060 = data_d1[239:232];
        6'd31: vec_data_060 = data_d1[247:240];
        6'd32: vec_data_060 = data_d1[255:248];
        6'd33: vec_data_060 = data_d1[263:256];
        6'd34: vec_data_060 = data_d1[271:264];
        6'd35: vec_data_060 = data_d1[279:272];
        6'd36: vec_data_060 = data_d1[287:280];
        6'd37: vec_data_060 = data_d1[295:288];
        6'd38: vec_data_060 = data_d1[303:296];
        6'd39: vec_data_060 = data_d1[311:304];
        6'd40: vec_data_060 = data_d1[319:312];
        6'd41: vec_data_060 = data_d1[327:320];
        6'd42: vec_data_060 = data_d1[335:328];
        6'd43: vec_data_060 = data_d1[343:336];
        6'd44: vec_data_060 = data_d1[351:344];
        6'd45: vec_data_060 = data_d1[359:352];
        6'd46: vec_data_060 = data_d1[367:360];
        6'd47: vec_data_060 = data_d1[375:368];
        6'd48: vec_data_060 = data_d1[383:376];
        6'd49: vec_data_060 = data_d1[391:384];
        6'd50: vec_data_060 = data_d1[399:392];
        6'd51: vec_data_060 = data_d1[407:400];
        6'd52: vec_data_060 = data_d1[415:408];
        6'd53: vec_data_060 = data_d1[423:416];
        6'd54: vec_data_060 = data_d1[431:424];
        6'd55: vec_data_060 = data_d1[439:432];
        6'd56: vec_data_060 = data_d1[447:440];
        6'd57: vec_data_060 = data_d1[455:448];
        6'd58: vec_data_060 = data_d1[463:456];
        6'd59: vec_data_060 = data_d1[471:464];
        6'd60: vec_data_060 = data_d1[479:472];
        6'd61: vec_data_060 = data_d1[487:480];
    endcase
end

always @(
  vec_sum_061_d1
  or data_d1
  ) begin
    vec_data_061 = 8'b0;
    case(vec_sum_061_d1)
        6'd1: vec_data_061 = data_d1[7:0];
        6'd2: vec_data_061 = data_d1[15:8];
        6'd3: vec_data_061 = data_d1[23:16];
        6'd4: vec_data_061 = data_d1[31:24];
        6'd5: vec_data_061 = data_d1[39:32];
        6'd6: vec_data_061 = data_d1[47:40];
        6'd7: vec_data_061 = data_d1[55:48];
        6'd8: vec_data_061 = data_d1[63:56];
        6'd9: vec_data_061 = data_d1[71:64];
        6'd10: vec_data_061 = data_d1[79:72];
        6'd11: vec_data_061 = data_d1[87:80];
        6'd12: vec_data_061 = data_d1[95:88];
        6'd13: vec_data_061 = data_d1[103:96];
        6'd14: vec_data_061 = data_d1[111:104];
        6'd15: vec_data_061 = data_d1[119:112];
        6'd16: vec_data_061 = data_d1[127:120];
        6'd17: vec_data_061 = data_d1[135:128];
        6'd18: vec_data_061 = data_d1[143:136];
        6'd19: vec_data_061 = data_d1[151:144];
        6'd20: vec_data_061 = data_d1[159:152];
        6'd21: vec_data_061 = data_d1[167:160];
        6'd22: vec_data_061 = data_d1[175:168];
        6'd23: vec_data_061 = data_d1[183:176];
        6'd24: vec_data_061 = data_d1[191:184];
        6'd25: vec_data_061 = data_d1[199:192];
        6'd26: vec_data_061 = data_d1[207:200];
        6'd27: vec_data_061 = data_d1[215:208];
        6'd28: vec_data_061 = data_d1[223:216];
        6'd29: vec_data_061 = data_d1[231:224];
        6'd30: vec_data_061 = data_d1[239:232];
        6'd31: vec_data_061 = data_d1[247:240];
        6'd32: vec_data_061 = data_d1[255:248];
        6'd33: vec_data_061 = data_d1[263:256];
        6'd34: vec_data_061 = data_d1[271:264];
        6'd35: vec_data_061 = data_d1[279:272];
        6'd36: vec_data_061 = data_d1[287:280];
        6'd37: vec_data_061 = data_d1[295:288];
        6'd38: vec_data_061 = data_d1[303:296];
        6'd39: vec_data_061 = data_d1[311:304];
        6'd40: vec_data_061 = data_d1[319:312];
        6'd41: vec_data_061 = data_d1[327:320];
        6'd42: vec_data_061 = data_d1[335:328];
        6'd43: vec_data_061 = data_d1[343:336];
        6'd44: vec_data_061 = data_d1[351:344];
        6'd45: vec_data_061 = data_d1[359:352];
        6'd46: vec_data_061 = data_d1[367:360];
        6'd47: vec_data_061 = data_d1[375:368];
        6'd48: vec_data_061 = data_d1[383:376];
        6'd49: vec_data_061 = data_d1[391:384];
        6'd50: vec_data_061 = data_d1[399:392];
        6'd51: vec_data_061 = data_d1[407:400];
        6'd52: vec_data_061 = data_d1[415:408];
        6'd53: vec_data_061 = data_d1[423:416];
        6'd54: vec_data_061 = data_d1[431:424];
        6'd55: vec_data_061 = data_d1[439:432];
        6'd56: vec_data_061 = data_d1[447:440];
        6'd57: vec_data_061 = data_d1[455:448];
        6'd58: vec_data_061 = data_d1[463:456];
        6'd59: vec_data_061 = data_d1[471:464];
        6'd60: vec_data_061 = data_d1[479:472];
        6'd61: vec_data_061 = data_d1[487:480];
        6'd62: vec_data_061 = data_d1[495:488];
    endcase
end

always @(
  vec_sum_062_d1
  or data_d1
  ) begin
    vec_data_062 = 8'b0;
    case(vec_sum_062_d1)
        6'd1: vec_data_062 = data_d1[7:0];
        6'd2: vec_data_062 = data_d1[15:8];
        6'd3: vec_data_062 = data_d1[23:16];
        6'd4: vec_data_062 = data_d1[31:24];
        6'd5: vec_data_062 = data_d1[39:32];
        6'd6: vec_data_062 = data_d1[47:40];
        6'd7: vec_data_062 = data_d1[55:48];
        6'd8: vec_data_062 = data_d1[63:56];
        6'd9: vec_data_062 = data_d1[71:64];
        6'd10: vec_data_062 = data_d1[79:72];
        6'd11: vec_data_062 = data_d1[87:80];
        6'd12: vec_data_062 = data_d1[95:88];
        6'd13: vec_data_062 = data_d1[103:96];
        6'd14: vec_data_062 = data_d1[111:104];
        6'd15: vec_data_062 = data_d1[119:112];
        6'd16: vec_data_062 = data_d1[127:120];
        6'd17: vec_data_062 = data_d1[135:128];
        6'd18: vec_data_062 = data_d1[143:136];
        6'd19: vec_data_062 = data_d1[151:144];
        6'd20: vec_data_062 = data_d1[159:152];
        6'd21: vec_data_062 = data_d1[167:160];
        6'd22: vec_data_062 = data_d1[175:168];
        6'd23: vec_data_062 = data_d1[183:176];
        6'd24: vec_data_062 = data_d1[191:184];
        6'd25: vec_data_062 = data_d1[199:192];
        6'd26: vec_data_062 = data_d1[207:200];
        6'd27: vec_data_062 = data_d1[215:208];
        6'd28: vec_data_062 = data_d1[223:216];
        6'd29: vec_data_062 = data_d1[231:224];
        6'd30: vec_data_062 = data_d1[239:232];
        6'd31: vec_data_062 = data_d1[247:240];
        6'd32: vec_data_062 = data_d1[255:248];
        6'd33: vec_data_062 = data_d1[263:256];
        6'd34: vec_data_062 = data_d1[271:264];
        6'd35: vec_data_062 = data_d1[279:272];
        6'd36: vec_data_062 = data_d1[287:280];
        6'd37: vec_data_062 = data_d1[295:288];
        6'd38: vec_data_062 = data_d1[303:296];
        6'd39: vec_data_062 = data_d1[311:304];
        6'd40: vec_data_062 = data_d1[319:312];
        6'd41: vec_data_062 = data_d1[327:320];
        6'd42: vec_data_062 = data_d1[335:328];
        6'd43: vec_data_062 = data_d1[343:336];
        6'd44: vec_data_062 = data_d1[351:344];
        6'd45: vec_data_062 = data_d1[359:352];
        6'd46: vec_data_062 = data_d1[367:360];
        6'd47: vec_data_062 = data_d1[375:368];
        6'd48: vec_data_062 = data_d1[383:376];
        6'd49: vec_data_062 = data_d1[391:384];
        6'd50: vec_data_062 = data_d1[399:392];
        6'd51: vec_data_062 = data_d1[407:400];
        6'd52: vec_data_062 = data_d1[415:408];
        6'd53: vec_data_062 = data_d1[423:416];
        6'd54: vec_data_062 = data_d1[431:424];
        6'd55: vec_data_062 = data_d1[439:432];
        6'd56: vec_data_062 = data_d1[447:440];
        6'd57: vec_data_062 = data_d1[455:448];
        6'd58: vec_data_062 = data_d1[463:456];
        6'd59: vec_data_062 = data_d1[471:464];
        6'd60: vec_data_062 = data_d1[479:472];
        6'd61: vec_data_062 = data_d1[487:480];
        6'd62: vec_data_062 = data_d1[495:488];
        6'd63: vec_data_062 = data_d1[503:496];
    endcase
end

always @(
  vec_sum_063_d1
  or data_d1
  ) begin
    vec_data_063 = 8'b0;
    case(vec_sum_063_d1)
        7'd1: vec_data_063 = data_d1[7:0];
        7'd2: vec_data_063 = data_d1[15:8];
        7'd3: vec_data_063 = data_d1[23:16];
        7'd4: vec_data_063 = data_d1[31:24];
        7'd5: vec_data_063 = data_d1[39:32];
        7'd6: vec_data_063 = data_d1[47:40];
        7'd7: vec_data_063 = data_d1[55:48];
        7'd8: vec_data_063 = data_d1[63:56];
        7'd9: vec_data_063 = data_d1[71:64];
        7'd10: vec_data_063 = data_d1[79:72];
        7'd11: vec_data_063 = data_d1[87:80];
        7'd12: vec_data_063 = data_d1[95:88];
        7'd13: vec_data_063 = data_d1[103:96];
        7'd14: vec_data_063 = data_d1[111:104];
        7'd15: vec_data_063 = data_d1[119:112];
        7'd16: vec_data_063 = data_d1[127:120];
        7'd17: vec_data_063 = data_d1[135:128];
        7'd18: vec_data_063 = data_d1[143:136];
        7'd19: vec_data_063 = data_d1[151:144];
        7'd20: vec_data_063 = data_d1[159:152];
        7'd21: vec_data_063 = data_d1[167:160];
        7'd22: vec_data_063 = data_d1[175:168];
        7'd23: vec_data_063 = data_d1[183:176];
        7'd24: vec_data_063 = data_d1[191:184];
        7'd25: vec_data_063 = data_d1[199:192];
        7'd26: vec_data_063 = data_d1[207:200];
        7'd27: vec_data_063 = data_d1[215:208];
        7'd28: vec_data_063 = data_d1[223:216];
        7'd29: vec_data_063 = data_d1[231:224];
        7'd30: vec_data_063 = data_d1[239:232];
        7'd31: vec_data_063 = data_d1[247:240];
        7'd32: vec_data_063 = data_d1[255:248];
        7'd33: vec_data_063 = data_d1[263:256];
        7'd34: vec_data_063 = data_d1[271:264];
        7'd35: vec_data_063 = data_d1[279:272];
        7'd36: vec_data_063 = data_d1[287:280];
        7'd37: vec_data_063 = data_d1[295:288];
        7'd38: vec_data_063 = data_d1[303:296];
        7'd39: vec_data_063 = data_d1[311:304];
        7'd40: vec_data_063 = data_d1[319:312];
        7'd41: vec_data_063 = data_d1[327:320];
        7'd42: vec_data_063 = data_d1[335:328];
        7'd43: vec_data_063 = data_d1[343:336];
        7'd44: vec_data_063 = data_d1[351:344];
        7'd45: vec_data_063 = data_d1[359:352];
        7'd46: vec_data_063 = data_d1[367:360];
        7'd47: vec_data_063 = data_d1[375:368];
        7'd48: vec_data_063 = data_d1[383:376];
        7'd49: vec_data_063 = data_d1[391:384];
        7'd50: vec_data_063 = data_d1[399:392];
        7'd51: vec_data_063 = data_d1[407:400];
        7'd52: vec_data_063 = data_d1[415:408];
        7'd53: vec_data_063 = data_d1[423:416];
        7'd54: vec_data_063 = data_d1[431:424];
        7'd55: vec_data_063 = data_d1[439:432];
        7'd56: vec_data_063 = data_d1[447:440];
        7'd57: vec_data_063 = data_d1[455:448];
        7'd58: vec_data_063 = data_d1[463:456];
        7'd59: vec_data_063 = data_d1[471:464];
        7'd60: vec_data_063 = data_d1[479:472];
        7'd61: vec_data_063 = data_d1[487:480];
        7'd62: vec_data_063 = data_d1[495:488];
        7'd63: vec_data_063 = data_d1[503:496];
        7'd64: vec_data_063 = data_d1[511:504];
    endcase
end

always @(
  vec_sum_064_d1
  or data_d1
  ) begin
    vec_data_064 = 8'b0;
    case(vec_sum_064_d1)
        7'd1: vec_data_064 = data_d1[7:0];
        7'd2: vec_data_064 = data_d1[15:8];
        7'd3: vec_data_064 = data_d1[23:16];
        7'd4: vec_data_064 = data_d1[31:24];
        7'd5: vec_data_064 = data_d1[39:32];
        7'd6: vec_data_064 = data_d1[47:40];
        7'd7: vec_data_064 = data_d1[55:48];
        7'd8: vec_data_064 = data_d1[63:56];
        7'd9: vec_data_064 = data_d1[71:64];
        7'd10: vec_data_064 = data_d1[79:72];
        7'd11: vec_data_064 = data_d1[87:80];
        7'd12: vec_data_064 = data_d1[95:88];
        7'd13: vec_data_064 = data_d1[103:96];
        7'd14: vec_data_064 = data_d1[111:104];
        7'd15: vec_data_064 = data_d1[119:112];
        7'd16: vec_data_064 = data_d1[127:120];
        7'd17: vec_data_064 = data_d1[135:128];
        7'd18: vec_data_064 = data_d1[143:136];
        7'd19: vec_data_064 = data_d1[151:144];
        7'd20: vec_data_064 = data_d1[159:152];
        7'd21: vec_data_064 = data_d1[167:160];
        7'd22: vec_data_064 = data_d1[175:168];
        7'd23: vec_data_064 = data_d1[183:176];
        7'd24: vec_data_064 = data_d1[191:184];
        7'd25: vec_data_064 = data_d1[199:192];
        7'd26: vec_data_064 = data_d1[207:200];
        7'd27: vec_data_064 = data_d1[215:208];
        7'd28: vec_data_064 = data_d1[223:216];
        7'd29: vec_data_064 = data_d1[231:224];
        7'd30: vec_data_064 = data_d1[239:232];
        7'd31: vec_data_064 = data_d1[247:240];
        7'd32: vec_data_064 = data_d1[255:248];
        7'd33: vec_data_064 = data_d1[263:256];
        7'd34: vec_data_064 = data_d1[271:264];
        7'd35: vec_data_064 = data_d1[279:272];
        7'd36: vec_data_064 = data_d1[287:280];
        7'd37: vec_data_064 = data_d1[295:288];
        7'd38: vec_data_064 = data_d1[303:296];
        7'd39: vec_data_064 = data_d1[311:304];
        7'd40: vec_data_064 = data_d1[319:312];
        7'd41: vec_data_064 = data_d1[327:320];
        7'd42: vec_data_064 = data_d1[335:328];
        7'd43: vec_data_064 = data_d1[343:336];
        7'd44: vec_data_064 = data_d1[351:344];
        7'd45: vec_data_064 = data_d1[359:352];
        7'd46: vec_data_064 = data_d1[367:360];
        7'd47: vec_data_064 = data_d1[375:368];
        7'd48: vec_data_064 = data_d1[383:376];
        7'd49: vec_data_064 = data_d1[391:384];
        7'd50: vec_data_064 = data_d1[399:392];
        7'd51: vec_data_064 = data_d1[407:400];
        7'd52: vec_data_064 = data_d1[415:408];
        7'd53: vec_data_064 = data_d1[423:416];
        7'd54: vec_data_064 = data_d1[431:424];
        7'd55: vec_data_064 = data_d1[439:432];
        7'd56: vec_data_064 = data_d1[447:440];
        7'd57: vec_data_064 = data_d1[455:448];
        7'd58: vec_data_064 = data_d1[463:456];
        7'd59: vec_data_064 = data_d1[471:464];
        7'd60: vec_data_064 = data_d1[479:472];
        7'd61: vec_data_064 = data_d1[487:480];
        7'd62: vec_data_064 = data_d1[495:488];
        7'd63: vec_data_064 = data_d1[503:496];
        7'd64: vec_data_064 = data_d1[511:504];
        7'd65: vec_data_064 = data_d1[519:512];
    endcase
end

always @(
  vec_sum_065_d1
  or data_d1
  ) begin
    vec_data_065 = 8'b0;
    case(vec_sum_065_d1)
        7'd1: vec_data_065 = data_d1[7:0];
        7'd2: vec_data_065 = data_d1[15:8];
        7'd3: vec_data_065 = data_d1[23:16];
        7'd4: vec_data_065 = data_d1[31:24];
        7'd5: vec_data_065 = data_d1[39:32];
        7'd6: vec_data_065 = data_d1[47:40];
        7'd7: vec_data_065 = data_d1[55:48];
        7'd8: vec_data_065 = data_d1[63:56];
        7'd9: vec_data_065 = data_d1[71:64];
        7'd10: vec_data_065 = data_d1[79:72];
        7'd11: vec_data_065 = data_d1[87:80];
        7'd12: vec_data_065 = data_d1[95:88];
        7'd13: vec_data_065 = data_d1[103:96];
        7'd14: vec_data_065 = data_d1[111:104];
        7'd15: vec_data_065 = data_d1[119:112];
        7'd16: vec_data_065 = data_d1[127:120];
        7'd17: vec_data_065 = data_d1[135:128];
        7'd18: vec_data_065 = data_d1[143:136];
        7'd19: vec_data_065 = data_d1[151:144];
        7'd20: vec_data_065 = data_d1[159:152];
        7'd21: vec_data_065 = data_d1[167:160];
        7'd22: vec_data_065 = data_d1[175:168];
        7'd23: vec_data_065 = data_d1[183:176];
        7'd24: vec_data_065 = data_d1[191:184];
        7'd25: vec_data_065 = data_d1[199:192];
        7'd26: vec_data_065 = data_d1[207:200];
        7'd27: vec_data_065 = data_d1[215:208];
        7'd28: vec_data_065 = data_d1[223:216];
        7'd29: vec_data_065 = data_d1[231:224];
        7'd30: vec_data_065 = data_d1[239:232];
        7'd31: vec_data_065 = data_d1[247:240];
        7'd32: vec_data_065 = data_d1[255:248];
        7'd33: vec_data_065 = data_d1[263:256];
        7'd34: vec_data_065 = data_d1[271:264];
        7'd35: vec_data_065 = data_d1[279:272];
        7'd36: vec_data_065 = data_d1[287:280];
        7'd37: vec_data_065 = data_d1[295:288];
        7'd38: vec_data_065 = data_d1[303:296];
        7'd39: vec_data_065 = data_d1[311:304];
        7'd40: vec_data_065 = data_d1[319:312];
        7'd41: vec_data_065 = data_d1[327:320];
        7'd42: vec_data_065 = data_d1[335:328];
        7'd43: vec_data_065 = data_d1[343:336];
        7'd44: vec_data_065 = data_d1[351:344];
        7'd45: vec_data_065 = data_d1[359:352];
        7'd46: vec_data_065 = data_d1[367:360];
        7'd47: vec_data_065 = data_d1[375:368];
        7'd48: vec_data_065 = data_d1[383:376];
        7'd49: vec_data_065 = data_d1[391:384];
        7'd50: vec_data_065 = data_d1[399:392];
        7'd51: vec_data_065 = data_d1[407:400];
        7'd52: vec_data_065 = data_d1[415:408];
        7'd53: vec_data_065 = data_d1[423:416];
        7'd54: vec_data_065 = data_d1[431:424];
        7'd55: vec_data_065 = data_d1[439:432];
        7'd56: vec_data_065 = data_d1[447:440];
        7'd57: vec_data_065 = data_d1[455:448];
        7'd58: vec_data_065 = data_d1[463:456];
        7'd59: vec_data_065 = data_d1[471:464];
        7'd60: vec_data_065 = data_d1[479:472];
        7'd61: vec_data_065 = data_d1[487:480];
        7'd62: vec_data_065 = data_d1[495:488];
        7'd63: vec_data_065 = data_d1[503:496];
        7'd64: vec_data_065 = data_d1[511:504];
        7'd65: vec_data_065 = data_d1[519:512];
        7'd66: vec_data_065 = data_d1[527:520];
    endcase
end

always @(
  vec_sum_066_d1
  or data_d1
  ) begin
    vec_data_066 = 8'b0;
    case(vec_sum_066_d1)
        7'd1: vec_data_066 = data_d1[7:0];
        7'd2: vec_data_066 = data_d1[15:8];
        7'd3: vec_data_066 = data_d1[23:16];
        7'd4: vec_data_066 = data_d1[31:24];
        7'd5: vec_data_066 = data_d1[39:32];
        7'd6: vec_data_066 = data_d1[47:40];
        7'd7: vec_data_066 = data_d1[55:48];
        7'd8: vec_data_066 = data_d1[63:56];
        7'd9: vec_data_066 = data_d1[71:64];
        7'd10: vec_data_066 = data_d1[79:72];
        7'd11: vec_data_066 = data_d1[87:80];
        7'd12: vec_data_066 = data_d1[95:88];
        7'd13: vec_data_066 = data_d1[103:96];
        7'd14: vec_data_066 = data_d1[111:104];
        7'd15: vec_data_066 = data_d1[119:112];
        7'd16: vec_data_066 = data_d1[127:120];
        7'd17: vec_data_066 = data_d1[135:128];
        7'd18: vec_data_066 = data_d1[143:136];
        7'd19: vec_data_066 = data_d1[151:144];
        7'd20: vec_data_066 = data_d1[159:152];
        7'd21: vec_data_066 = data_d1[167:160];
        7'd22: vec_data_066 = data_d1[175:168];
        7'd23: vec_data_066 = data_d1[183:176];
        7'd24: vec_data_066 = data_d1[191:184];
        7'd25: vec_data_066 = data_d1[199:192];
        7'd26: vec_data_066 = data_d1[207:200];
        7'd27: vec_data_066 = data_d1[215:208];
        7'd28: vec_data_066 = data_d1[223:216];
        7'd29: vec_data_066 = data_d1[231:224];
        7'd30: vec_data_066 = data_d1[239:232];
        7'd31: vec_data_066 = data_d1[247:240];
        7'd32: vec_data_066 = data_d1[255:248];
        7'd33: vec_data_066 = data_d1[263:256];
        7'd34: vec_data_066 = data_d1[271:264];
        7'd35: vec_data_066 = data_d1[279:272];
        7'd36: vec_data_066 = data_d1[287:280];
        7'd37: vec_data_066 = data_d1[295:288];
        7'd38: vec_data_066 = data_d1[303:296];
        7'd39: vec_data_066 = data_d1[311:304];
        7'd40: vec_data_066 = data_d1[319:312];
        7'd41: vec_data_066 = data_d1[327:320];
        7'd42: vec_data_066 = data_d1[335:328];
        7'd43: vec_data_066 = data_d1[343:336];
        7'd44: vec_data_066 = data_d1[351:344];
        7'd45: vec_data_066 = data_d1[359:352];
        7'd46: vec_data_066 = data_d1[367:360];
        7'd47: vec_data_066 = data_d1[375:368];
        7'd48: vec_data_066 = data_d1[383:376];
        7'd49: vec_data_066 = data_d1[391:384];
        7'd50: vec_data_066 = data_d1[399:392];
        7'd51: vec_data_066 = data_d1[407:400];
        7'd52: vec_data_066 = data_d1[415:408];
        7'd53: vec_data_066 = data_d1[423:416];
        7'd54: vec_data_066 = data_d1[431:424];
        7'd55: vec_data_066 = data_d1[439:432];
        7'd56: vec_data_066 = data_d1[447:440];
        7'd57: vec_data_066 = data_d1[455:448];
        7'd58: vec_data_066 = data_d1[463:456];
        7'd59: vec_data_066 = data_d1[471:464];
        7'd60: vec_data_066 = data_d1[479:472];
        7'd61: vec_data_066 = data_d1[487:480];
        7'd62: vec_data_066 = data_d1[495:488];
        7'd63: vec_data_066 = data_d1[503:496];
        7'd64: vec_data_066 = data_d1[511:504];
        7'd65: vec_data_066 = data_d1[519:512];
        7'd66: vec_data_066 = data_d1[527:520];
        7'd67: vec_data_066 = data_d1[535:528];
    endcase
end

always @(
  vec_sum_067_d1
  or data_d1
  ) begin
    vec_data_067 = 8'b0;
    case(vec_sum_067_d1)
        7'd1: vec_data_067 = data_d1[7:0];
        7'd2: vec_data_067 = data_d1[15:8];
        7'd3: vec_data_067 = data_d1[23:16];
        7'd4: vec_data_067 = data_d1[31:24];
        7'd5: vec_data_067 = data_d1[39:32];
        7'd6: vec_data_067 = data_d1[47:40];
        7'd7: vec_data_067 = data_d1[55:48];
        7'd8: vec_data_067 = data_d1[63:56];
        7'd9: vec_data_067 = data_d1[71:64];
        7'd10: vec_data_067 = data_d1[79:72];
        7'd11: vec_data_067 = data_d1[87:80];
        7'd12: vec_data_067 = data_d1[95:88];
        7'd13: vec_data_067 = data_d1[103:96];
        7'd14: vec_data_067 = data_d1[111:104];
        7'd15: vec_data_067 = data_d1[119:112];
        7'd16: vec_data_067 = data_d1[127:120];
        7'd17: vec_data_067 = data_d1[135:128];
        7'd18: vec_data_067 = data_d1[143:136];
        7'd19: vec_data_067 = data_d1[151:144];
        7'd20: vec_data_067 = data_d1[159:152];
        7'd21: vec_data_067 = data_d1[167:160];
        7'd22: vec_data_067 = data_d1[175:168];
        7'd23: vec_data_067 = data_d1[183:176];
        7'd24: vec_data_067 = data_d1[191:184];
        7'd25: vec_data_067 = data_d1[199:192];
        7'd26: vec_data_067 = data_d1[207:200];
        7'd27: vec_data_067 = data_d1[215:208];
        7'd28: vec_data_067 = data_d1[223:216];
        7'd29: vec_data_067 = data_d1[231:224];
        7'd30: vec_data_067 = data_d1[239:232];
        7'd31: vec_data_067 = data_d1[247:240];
        7'd32: vec_data_067 = data_d1[255:248];
        7'd33: vec_data_067 = data_d1[263:256];
        7'd34: vec_data_067 = data_d1[271:264];
        7'd35: vec_data_067 = data_d1[279:272];
        7'd36: vec_data_067 = data_d1[287:280];
        7'd37: vec_data_067 = data_d1[295:288];
        7'd38: vec_data_067 = data_d1[303:296];
        7'd39: vec_data_067 = data_d1[311:304];
        7'd40: vec_data_067 = data_d1[319:312];
        7'd41: vec_data_067 = data_d1[327:320];
        7'd42: vec_data_067 = data_d1[335:328];
        7'd43: vec_data_067 = data_d1[343:336];
        7'd44: vec_data_067 = data_d1[351:344];
        7'd45: vec_data_067 = data_d1[359:352];
        7'd46: vec_data_067 = data_d1[367:360];
        7'd47: vec_data_067 = data_d1[375:368];
        7'd48: vec_data_067 = data_d1[383:376];
        7'd49: vec_data_067 = data_d1[391:384];
        7'd50: vec_data_067 = data_d1[399:392];
        7'd51: vec_data_067 = data_d1[407:400];
        7'd52: vec_data_067 = data_d1[415:408];
        7'd53: vec_data_067 = data_d1[423:416];
        7'd54: vec_data_067 = data_d1[431:424];
        7'd55: vec_data_067 = data_d1[439:432];
        7'd56: vec_data_067 = data_d1[447:440];
        7'd57: vec_data_067 = data_d1[455:448];
        7'd58: vec_data_067 = data_d1[463:456];
        7'd59: vec_data_067 = data_d1[471:464];
        7'd60: vec_data_067 = data_d1[479:472];
        7'd61: vec_data_067 = data_d1[487:480];
        7'd62: vec_data_067 = data_d1[495:488];
        7'd63: vec_data_067 = data_d1[503:496];
        7'd64: vec_data_067 = data_d1[511:504];
        7'd65: vec_data_067 = data_d1[519:512];
        7'd66: vec_data_067 = data_d1[527:520];
        7'd67: vec_data_067 = data_d1[535:528];
        7'd68: vec_data_067 = data_d1[543:536];
    endcase
end

always @(
  vec_sum_068_d1
  or data_d1
  ) begin
    vec_data_068 = 8'b0;
    case(vec_sum_068_d1)
        7'd1: vec_data_068 = data_d1[7:0];
        7'd2: vec_data_068 = data_d1[15:8];
        7'd3: vec_data_068 = data_d1[23:16];
        7'd4: vec_data_068 = data_d1[31:24];
        7'd5: vec_data_068 = data_d1[39:32];
        7'd6: vec_data_068 = data_d1[47:40];
        7'd7: vec_data_068 = data_d1[55:48];
        7'd8: vec_data_068 = data_d1[63:56];
        7'd9: vec_data_068 = data_d1[71:64];
        7'd10: vec_data_068 = data_d1[79:72];
        7'd11: vec_data_068 = data_d1[87:80];
        7'd12: vec_data_068 = data_d1[95:88];
        7'd13: vec_data_068 = data_d1[103:96];
        7'd14: vec_data_068 = data_d1[111:104];
        7'd15: vec_data_068 = data_d1[119:112];
        7'd16: vec_data_068 = data_d1[127:120];
        7'd17: vec_data_068 = data_d1[135:128];
        7'd18: vec_data_068 = data_d1[143:136];
        7'd19: vec_data_068 = data_d1[151:144];
        7'd20: vec_data_068 = data_d1[159:152];
        7'd21: vec_data_068 = data_d1[167:160];
        7'd22: vec_data_068 = data_d1[175:168];
        7'd23: vec_data_068 = data_d1[183:176];
        7'd24: vec_data_068 = data_d1[191:184];
        7'd25: vec_data_068 = data_d1[199:192];
        7'd26: vec_data_068 = data_d1[207:200];
        7'd27: vec_data_068 = data_d1[215:208];
        7'd28: vec_data_068 = data_d1[223:216];
        7'd29: vec_data_068 = data_d1[231:224];
        7'd30: vec_data_068 = data_d1[239:232];
        7'd31: vec_data_068 = data_d1[247:240];
        7'd32: vec_data_068 = data_d1[255:248];
        7'd33: vec_data_068 = data_d1[263:256];
        7'd34: vec_data_068 = data_d1[271:264];
        7'd35: vec_data_068 = data_d1[279:272];
        7'd36: vec_data_068 = data_d1[287:280];
        7'd37: vec_data_068 = data_d1[295:288];
        7'd38: vec_data_068 = data_d1[303:296];
        7'd39: vec_data_068 = data_d1[311:304];
        7'd40: vec_data_068 = data_d1[319:312];
        7'd41: vec_data_068 = data_d1[327:320];
        7'd42: vec_data_068 = data_d1[335:328];
        7'd43: vec_data_068 = data_d1[343:336];
        7'd44: vec_data_068 = data_d1[351:344];
        7'd45: vec_data_068 = data_d1[359:352];
        7'd46: vec_data_068 = data_d1[367:360];
        7'd47: vec_data_068 = data_d1[375:368];
        7'd48: vec_data_068 = data_d1[383:376];
        7'd49: vec_data_068 = data_d1[391:384];
        7'd50: vec_data_068 = data_d1[399:392];
        7'd51: vec_data_068 = data_d1[407:400];
        7'd52: vec_data_068 = data_d1[415:408];
        7'd53: vec_data_068 = data_d1[423:416];
        7'd54: vec_data_068 = data_d1[431:424];
        7'd55: vec_data_068 = data_d1[439:432];
        7'd56: vec_data_068 = data_d1[447:440];
        7'd57: vec_data_068 = data_d1[455:448];
        7'd58: vec_data_068 = data_d1[463:456];
        7'd59: vec_data_068 = data_d1[471:464];
        7'd60: vec_data_068 = data_d1[479:472];
        7'd61: vec_data_068 = data_d1[487:480];
        7'd62: vec_data_068 = data_d1[495:488];
        7'd63: vec_data_068 = data_d1[503:496];
        7'd64: vec_data_068 = data_d1[511:504];
        7'd65: vec_data_068 = data_d1[519:512];
        7'd66: vec_data_068 = data_d1[527:520];
        7'd67: vec_data_068 = data_d1[535:528];
        7'd68: vec_data_068 = data_d1[543:536];
        7'd69: vec_data_068 = data_d1[551:544];
    endcase
end

always @(
  vec_sum_069_d1
  or data_d1
  ) begin
    vec_data_069 = 8'b0;
    case(vec_sum_069_d1)
        7'd1: vec_data_069 = data_d1[7:0];
        7'd2: vec_data_069 = data_d1[15:8];
        7'd3: vec_data_069 = data_d1[23:16];
        7'd4: vec_data_069 = data_d1[31:24];
        7'd5: vec_data_069 = data_d1[39:32];
        7'd6: vec_data_069 = data_d1[47:40];
        7'd7: vec_data_069 = data_d1[55:48];
        7'd8: vec_data_069 = data_d1[63:56];
        7'd9: vec_data_069 = data_d1[71:64];
        7'd10: vec_data_069 = data_d1[79:72];
        7'd11: vec_data_069 = data_d1[87:80];
        7'd12: vec_data_069 = data_d1[95:88];
        7'd13: vec_data_069 = data_d1[103:96];
        7'd14: vec_data_069 = data_d1[111:104];
        7'd15: vec_data_069 = data_d1[119:112];
        7'd16: vec_data_069 = data_d1[127:120];
        7'd17: vec_data_069 = data_d1[135:128];
        7'd18: vec_data_069 = data_d1[143:136];
        7'd19: vec_data_069 = data_d1[151:144];
        7'd20: vec_data_069 = data_d1[159:152];
        7'd21: vec_data_069 = data_d1[167:160];
        7'd22: vec_data_069 = data_d1[175:168];
        7'd23: vec_data_069 = data_d1[183:176];
        7'd24: vec_data_069 = data_d1[191:184];
        7'd25: vec_data_069 = data_d1[199:192];
        7'd26: vec_data_069 = data_d1[207:200];
        7'd27: vec_data_069 = data_d1[215:208];
        7'd28: vec_data_069 = data_d1[223:216];
        7'd29: vec_data_069 = data_d1[231:224];
        7'd30: vec_data_069 = data_d1[239:232];
        7'd31: vec_data_069 = data_d1[247:240];
        7'd32: vec_data_069 = data_d1[255:248];
        7'd33: vec_data_069 = data_d1[263:256];
        7'd34: vec_data_069 = data_d1[271:264];
        7'd35: vec_data_069 = data_d1[279:272];
        7'd36: vec_data_069 = data_d1[287:280];
        7'd37: vec_data_069 = data_d1[295:288];
        7'd38: vec_data_069 = data_d1[303:296];
        7'd39: vec_data_069 = data_d1[311:304];
        7'd40: vec_data_069 = data_d1[319:312];
        7'd41: vec_data_069 = data_d1[327:320];
        7'd42: vec_data_069 = data_d1[335:328];
        7'd43: vec_data_069 = data_d1[343:336];
        7'd44: vec_data_069 = data_d1[351:344];
        7'd45: vec_data_069 = data_d1[359:352];
        7'd46: vec_data_069 = data_d1[367:360];
        7'd47: vec_data_069 = data_d1[375:368];
        7'd48: vec_data_069 = data_d1[383:376];
        7'd49: vec_data_069 = data_d1[391:384];
        7'd50: vec_data_069 = data_d1[399:392];
        7'd51: vec_data_069 = data_d1[407:400];
        7'd52: vec_data_069 = data_d1[415:408];
        7'd53: vec_data_069 = data_d1[423:416];
        7'd54: vec_data_069 = data_d1[431:424];
        7'd55: vec_data_069 = data_d1[439:432];
        7'd56: vec_data_069 = data_d1[447:440];
        7'd57: vec_data_069 = data_d1[455:448];
        7'd58: vec_data_069 = data_d1[463:456];
        7'd59: vec_data_069 = data_d1[471:464];
        7'd60: vec_data_069 = data_d1[479:472];
        7'd61: vec_data_069 = data_d1[487:480];
        7'd62: vec_data_069 = data_d1[495:488];
        7'd63: vec_data_069 = data_d1[503:496];
        7'd64: vec_data_069 = data_d1[511:504];
        7'd65: vec_data_069 = data_d1[519:512];
        7'd66: vec_data_069 = data_d1[527:520];
        7'd67: vec_data_069 = data_d1[535:528];
        7'd68: vec_data_069 = data_d1[543:536];
        7'd69: vec_data_069 = data_d1[551:544];
        7'd70: vec_data_069 = data_d1[559:552];
    endcase
end

always @(
  vec_sum_070_d1
  or data_d1
  ) begin
    vec_data_070 = 8'b0;
    case(vec_sum_070_d1)
        7'd1: vec_data_070 = data_d1[7:0];
        7'd2: vec_data_070 = data_d1[15:8];
        7'd3: vec_data_070 = data_d1[23:16];
        7'd4: vec_data_070 = data_d1[31:24];
        7'd5: vec_data_070 = data_d1[39:32];
        7'd6: vec_data_070 = data_d1[47:40];
        7'd7: vec_data_070 = data_d1[55:48];
        7'd8: vec_data_070 = data_d1[63:56];
        7'd9: vec_data_070 = data_d1[71:64];
        7'd10: vec_data_070 = data_d1[79:72];
        7'd11: vec_data_070 = data_d1[87:80];
        7'd12: vec_data_070 = data_d1[95:88];
        7'd13: vec_data_070 = data_d1[103:96];
        7'd14: vec_data_070 = data_d1[111:104];
        7'd15: vec_data_070 = data_d1[119:112];
        7'd16: vec_data_070 = data_d1[127:120];
        7'd17: vec_data_070 = data_d1[135:128];
        7'd18: vec_data_070 = data_d1[143:136];
        7'd19: vec_data_070 = data_d1[151:144];
        7'd20: vec_data_070 = data_d1[159:152];
        7'd21: vec_data_070 = data_d1[167:160];
        7'd22: vec_data_070 = data_d1[175:168];
        7'd23: vec_data_070 = data_d1[183:176];
        7'd24: vec_data_070 = data_d1[191:184];
        7'd25: vec_data_070 = data_d1[199:192];
        7'd26: vec_data_070 = data_d1[207:200];
        7'd27: vec_data_070 = data_d1[215:208];
        7'd28: vec_data_070 = data_d1[223:216];
        7'd29: vec_data_070 = data_d1[231:224];
        7'd30: vec_data_070 = data_d1[239:232];
        7'd31: vec_data_070 = data_d1[247:240];
        7'd32: vec_data_070 = data_d1[255:248];
        7'd33: vec_data_070 = data_d1[263:256];
        7'd34: vec_data_070 = data_d1[271:264];
        7'd35: vec_data_070 = data_d1[279:272];
        7'd36: vec_data_070 = data_d1[287:280];
        7'd37: vec_data_070 = data_d1[295:288];
        7'd38: vec_data_070 = data_d1[303:296];
        7'd39: vec_data_070 = data_d1[311:304];
        7'd40: vec_data_070 = data_d1[319:312];
        7'd41: vec_data_070 = data_d1[327:320];
        7'd42: vec_data_070 = data_d1[335:328];
        7'd43: vec_data_070 = data_d1[343:336];
        7'd44: vec_data_070 = data_d1[351:344];
        7'd45: vec_data_070 = data_d1[359:352];
        7'd46: vec_data_070 = data_d1[367:360];
        7'd47: vec_data_070 = data_d1[375:368];
        7'd48: vec_data_070 = data_d1[383:376];
        7'd49: vec_data_070 = data_d1[391:384];
        7'd50: vec_data_070 = data_d1[399:392];
        7'd51: vec_data_070 = data_d1[407:400];
        7'd52: vec_data_070 = data_d1[415:408];
        7'd53: vec_data_070 = data_d1[423:416];
        7'd54: vec_data_070 = data_d1[431:424];
        7'd55: vec_data_070 = data_d1[439:432];
        7'd56: vec_data_070 = data_d1[447:440];
        7'd57: vec_data_070 = data_d1[455:448];
        7'd58: vec_data_070 = data_d1[463:456];
        7'd59: vec_data_070 = data_d1[471:464];
        7'd60: vec_data_070 = data_d1[479:472];
        7'd61: vec_data_070 = data_d1[487:480];
        7'd62: vec_data_070 = data_d1[495:488];
        7'd63: vec_data_070 = data_d1[503:496];
        7'd64: vec_data_070 = data_d1[511:504];
        7'd65: vec_data_070 = data_d1[519:512];
        7'd66: vec_data_070 = data_d1[527:520];
        7'd67: vec_data_070 = data_d1[535:528];
        7'd68: vec_data_070 = data_d1[543:536];
        7'd69: vec_data_070 = data_d1[551:544];
        7'd70: vec_data_070 = data_d1[559:552];
        7'd71: vec_data_070 = data_d1[567:560];
    endcase
end

always @(
  vec_sum_071_d1
  or data_d1
  ) begin
    vec_data_071 = 8'b0;
    case(vec_sum_071_d1)
        7'd1: vec_data_071 = data_d1[7:0];
        7'd2: vec_data_071 = data_d1[15:8];
        7'd3: vec_data_071 = data_d1[23:16];
        7'd4: vec_data_071 = data_d1[31:24];
        7'd5: vec_data_071 = data_d1[39:32];
        7'd6: vec_data_071 = data_d1[47:40];
        7'd7: vec_data_071 = data_d1[55:48];
        7'd8: vec_data_071 = data_d1[63:56];
        7'd9: vec_data_071 = data_d1[71:64];
        7'd10: vec_data_071 = data_d1[79:72];
        7'd11: vec_data_071 = data_d1[87:80];
        7'd12: vec_data_071 = data_d1[95:88];
        7'd13: vec_data_071 = data_d1[103:96];
        7'd14: vec_data_071 = data_d1[111:104];
        7'd15: vec_data_071 = data_d1[119:112];
        7'd16: vec_data_071 = data_d1[127:120];
        7'd17: vec_data_071 = data_d1[135:128];
        7'd18: vec_data_071 = data_d1[143:136];
        7'd19: vec_data_071 = data_d1[151:144];
        7'd20: vec_data_071 = data_d1[159:152];
        7'd21: vec_data_071 = data_d1[167:160];
        7'd22: vec_data_071 = data_d1[175:168];
        7'd23: vec_data_071 = data_d1[183:176];
        7'd24: vec_data_071 = data_d1[191:184];
        7'd25: vec_data_071 = data_d1[199:192];
        7'd26: vec_data_071 = data_d1[207:200];
        7'd27: vec_data_071 = data_d1[215:208];
        7'd28: vec_data_071 = data_d1[223:216];
        7'd29: vec_data_071 = data_d1[231:224];
        7'd30: vec_data_071 = data_d1[239:232];
        7'd31: vec_data_071 = data_d1[247:240];
        7'd32: vec_data_071 = data_d1[255:248];
        7'd33: vec_data_071 = data_d1[263:256];
        7'd34: vec_data_071 = data_d1[271:264];
        7'd35: vec_data_071 = data_d1[279:272];
        7'd36: vec_data_071 = data_d1[287:280];
        7'd37: vec_data_071 = data_d1[295:288];
        7'd38: vec_data_071 = data_d1[303:296];
        7'd39: vec_data_071 = data_d1[311:304];
        7'd40: vec_data_071 = data_d1[319:312];
        7'd41: vec_data_071 = data_d1[327:320];
        7'd42: vec_data_071 = data_d1[335:328];
        7'd43: vec_data_071 = data_d1[343:336];
        7'd44: vec_data_071 = data_d1[351:344];
        7'd45: vec_data_071 = data_d1[359:352];
        7'd46: vec_data_071 = data_d1[367:360];
        7'd47: vec_data_071 = data_d1[375:368];
        7'd48: vec_data_071 = data_d1[383:376];
        7'd49: vec_data_071 = data_d1[391:384];
        7'd50: vec_data_071 = data_d1[399:392];
        7'd51: vec_data_071 = data_d1[407:400];
        7'd52: vec_data_071 = data_d1[415:408];
        7'd53: vec_data_071 = data_d1[423:416];
        7'd54: vec_data_071 = data_d1[431:424];
        7'd55: vec_data_071 = data_d1[439:432];
        7'd56: vec_data_071 = data_d1[447:440];
        7'd57: vec_data_071 = data_d1[455:448];
        7'd58: vec_data_071 = data_d1[463:456];
        7'd59: vec_data_071 = data_d1[471:464];
        7'd60: vec_data_071 = data_d1[479:472];
        7'd61: vec_data_071 = data_d1[487:480];
        7'd62: vec_data_071 = data_d1[495:488];
        7'd63: vec_data_071 = data_d1[503:496];
        7'd64: vec_data_071 = data_d1[511:504];
        7'd65: vec_data_071 = data_d1[519:512];
        7'd66: vec_data_071 = data_d1[527:520];
        7'd67: vec_data_071 = data_d1[535:528];
        7'd68: vec_data_071 = data_d1[543:536];
        7'd69: vec_data_071 = data_d1[551:544];
        7'd70: vec_data_071 = data_d1[559:552];
        7'd71: vec_data_071 = data_d1[567:560];
        7'd72: vec_data_071 = data_d1[575:568];
    endcase
end

always @(
  vec_sum_072_d1
  or data_d1
  ) begin
    vec_data_072 = 8'b0;
    case(vec_sum_072_d1)
        7'd1: vec_data_072 = data_d1[7:0];
        7'd2: vec_data_072 = data_d1[15:8];
        7'd3: vec_data_072 = data_d1[23:16];
        7'd4: vec_data_072 = data_d1[31:24];
        7'd5: vec_data_072 = data_d1[39:32];
        7'd6: vec_data_072 = data_d1[47:40];
        7'd7: vec_data_072 = data_d1[55:48];
        7'd8: vec_data_072 = data_d1[63:56];
        7'd9: vec_data_072 = data_d1[71:64];
        7'd10: vec_data_072 = data_d1[79:72];
        7'd11: vec_data_072 = data_d1[87:80];
        7'd12: vec_data_072 = data_d1[95:88];
        7'd13: vec_data_072 = data_d1[103:96];
        7'd14: vec_data_072 = data_d1[111:104];
        7'd15: vec_data_072 = data_d1[119:112];
        7'd16: vec_data_072 = data_d1[127:120];
        7'd17: vec_data_072 = data_d1[135:128];
        7'd18: vec_data_072 = data_d1[143:136];
        7'd19: vec_data_072 = data_d1[151:144];
        7'd20: vec_data_072 = data_d1[159:152];
        7'd21: vec_data_072 = data_d1[167:160];
        7'd22: vec_data_072 = data_d1[175:168];
        7'd23: vec_data_072 = data_d1[183:176];
        7'd24: vec_data_072 = data_d1[191:184];
        7'd25: vec_data_072 = data_d1[199:192];
        7'd26: vec_data_072 = data_d1[207:200];
        7'd27: vec_data_072 = data_d1[215:208];
        7'd28: vec_data_072 = data_d1[223:216];
        7'd29: vec_data_072 = data_d1[231:224];
        7'd30: vec_data_072 = data_d1[239:232];
        7'd31: vec_data_072 = data_d1[247:240];
        7'd32: vec_data_072 = data_d1[255:248];
        7'd33: vec_data_072 = data_d1[263:256];
        7'd34: vec_data_072 = data_d1[271:264];
        7'd35: vec_data_072 = data_d1[279:272];
        7'd36: vec_data_072 = data_d1[287:280];
        7'd37: vec_data_072 = data_d1[295:288];
        7'd38: vec_data_072 = data_d1[303:296];
        7'd39: vec_data_072 = data_d1[311:304];
        7'd40: vec_data_072 = data_d1[319:312];
        7'd41: vec_data_072 = data_d1[327:320];
        7'd42: vec_data_072 = data_d1[335:328];
        7'd43: vec_data_072 = data_d1[343:336];
        7'd44: vec_data_072 = data_d1[351:344];
        7'd45: vec_data_072 = data_d1[359:352];
        7'd46: vec_data_072 = data_d1[367:360];
        7'd47: vec_data_072 = data_d1[375:368];
        7'd48: vec_data_072 = data_d1[383:376];
        7'd49: vec_data_072 = data_d1[391:384];
        7'd50: vec_data_072 = data_d1[399:392];
        7'd51: vec_data_072 = data_d1[407:400];
        7'd52: vec_data_072 = data_d1[415:408];
        7'd53: vec_data_072 = data_d1[423:416];
        7'd54: vec_data_072 = data_d1[431:424];
        7'd55: vec_data_072 = data_d1[439:432];
        7'd56: vec_data_072 = data_d1[447:440];
        7'd57: vec_data_072 = data_d1[455:448];
        7'd58: vec_data_072 = data_d1[463:456];
        7'd59: vec_data_072 = data_d1[471:464];
        7'd60: vec_data_072 = data_d1[479:472];
        7'd61: vec_data_072 = data_d1[487:480];
        7'd62: vec_data_072 = data_d1[495:488];
        7'd63: vec_data_072 = data_d1[503:496];
        7'd64: vec_data_072 = data_d1[511:504];
        7'd65: vec_data_072 = data_d1[519:512];
        7'd66: vec_data_072 = data_d1[527:520];
        7'd67: vec_data_072 = data_d1[535:528];
        7'd68: vec_data_072 = data_d1[543:536];
        7'd69: vec_data_072 = data_d1[551:544];
        7'd70: vec_data_072 = data_d1[559:552];
        7'd71: vec_data_072 = data_d1[567:560];
        7'd72: vec_data_072 = data_d1[575:568];
        7'd73: vec_data_072 = data_d1[583:576];
    endcase
end

always @(
  vec_sum_073_d1
  or data_d1
  ) begin
    vec_data_073 = 8'b0;
    case(vec_sum_073_d1)
        7'd1: vec_data_073 = data_d1[7:0];
        7'd2: vec_data_073 = data_d1[15:8];
        7'd3: vec_data_073 = data_d1[23:16];
        7'd4: vec_data_073 = data_d1[31:24];
        7'd5: vec_data_073 = data_d1[39:32];
        7'd6: vec_data_073 = data_d1[47:40];
        7'd7: vec_data_073 = data_d1[55:48];
        7'd8: vec_data_073 = data_d1[63:56];
        7'd9: vec_data_073 = data_d1[71:64];
        7'd10: vec_data_073 = data_d1[79:72];
        7'd11: vec_data_073 = data_d1[87:80];
        7'd12: vec_data_073 = data_d1[95:88];
        7'd13: vec_data_073 = data_d1[103:96];
        7'd14: vec_data_073 = data_d1[111:104];
        7'd15: vec_data_073 = data_d1[119:112];
        7'd16: vec_data_073 = data_d1[127:120];
        7'd17: vec_data_073 = data_d1[135:128];
        7'd18: vec_data_073 = data_d1[143:136];
        7'd19: vec_data_073 = data_d1[151:144];
        7'd20: vec_data_073 = data_d1[159:152];
        7'd21: vec_data_073 = data_d1[167:160];
        7'd22: vec_data_073 = data_d1[175:168];
        7'd23: vec_data_073 = data_d1[183:176];
        7'd24: vec_data_073 = data_d1[191:184];
        7'd25: vec_data_073 = data_d1[199:192];
        7'd26: vec_data_073 = data_d1[207:200];
        7'd27: vec_data_073 = data_d1[215:208];
        7'd28: vec_data_073 = data_d1[223:216];
        7'd29: vec_data_073 = data_d1[231:224];
        7'd30: vec_data_073 = data_d1[239:232];
        7'd31: vec_data_073 = data_d1[247:240];
        7'd32: vec_data_073 = data_d1[255:248];
        7'd33: vec_data_073 = data_d1[263:256];
        7'd34: vec_data_073 = data_d1[271:264];
        7'd35: vec_data_073 = data_d1[279:272];
        7'd36: vec_data_073 = data_d1[287:280];
        7'd37: vec_data_073 = data_d1[295:288];
        7'd38: vec_data_073 = data_d1[303:296];
        7'd39: vec_data_073 = data_d1[311:304];
        7'd40: vec_data_073 = data_d1[319:312];
        7'd41: vec_data_073 = data_d1[327:320];
        7'd42: vec_data_073 = data_d1[335:328];
        7'd43: vec_data_073 = data_d1[343:336];
        7'd44: vec_data_073 = data_d1[351:344];
        7'd45: vec_data_073 = data_d1[359:352];
        7'd46: vec_data_073 = data_d1[367:360];
        7'd47: vec_data_073 = data_d1[375:368];
        7'd48: vec_data_073 = data_d1[383:376];
        7'd49: vec_data_073 = data_d1[391:384];
        7'd50: vec_data_073 = data_d1[399:392];
        7'd51: vec_data_073 = data_d1[407:400];
        7'd52: vec_data_073 = data_d1[415:408];
        7'd53: vec_data_073 = data_d1[423:416];
        7'd54: vec_data_073 = data_d1[431:424];
        7'd55: vec_data_073 = data_d1[439:432];
        7'd56: vec_data_073 = data_d1[447:440];
        7'd57: vec_data_073 = data_d1[455:448];
        7'd58: vec_data_073 = data_d1[463:456];
        7'd59: vec_data_073 = data_d1[471:464];
        7'd60: vec_data_073 = data_d1[479:472];
        7'd61: vec_data_073 = data_d1[487:480];
        7'd62: vec_data_073 = data_d1[495:488];
        7'd63: vec_data_073 = data_d1[503:496];
        7'd64: vec_data_073 = data_d1[511:504];
        7'd65: vec_data_073 = data_d1[519:512];
        7'd66: vec_data_073 = data_d1[527:520];
        7'd67: vec_data_073 = data_d1[535:528];
        7'd68: vec_data_073 = data_d1[543:536];
        7'd69: vec_data_073 = data_d1[551:544];
        7'd70: vec_data_073 = data_d1[559:552];
        7'd71: vec_data_073 = data_d1[567:560];
        7'd72: vec_data_073 = data_d1[575:568];
        7'd73: vec_data_073 = data_d1[583:576];
        7'd74: vec_data_073 = data_d1[591:584];
    endcase
end

always @(
  vec_sum_074_d1
  or data_d1
  ) begin
    vec_data_074 = 8'b0;
    case(vec_sum_074_d1)
        7'd1: vec_data_074 = data_d1[7:0];
        7'd2: vec_data_074 = data_d1[15:8];
        7'd3: vec_data_074 = data_d1[23:16];
        7'd4: vec_data_074 = data_d1[31:24];
        7'd5: vec_data_074 = data_d1[39:32];
        7'd6: vec_data_074 = data_d1[47:40];
        7'd7: vec_data_074 = data_d1[55:48];
        7'd8: vec_data_074 = data_d1[63:56];
        7'd9: vec_data_074 = data_d1[71:64];
        7'd10: vec_data_074 = data_d1[79:72];
        7'd11: vec_data_074 = data_d1[87:80];
        7'd12: vec_data_074 = data_d1[95:88];
        7'd13: vec_data_074 = data_d1[103:96];
        7'd14: vec_data_074 = data_d1[111:104];
        7'd15: vec_data_074 = data_d1[119:112];
        7'd16: vec_data_074 = data_d1[127:120];
        7'd17: vec_data_074 = data_d1[135:128];
        7'd18: vec_data_074 = data_d1[143:136];
        7'd19: vec_data_074 = data_d1[151:144];
        7'd20: vec_data_074 = data_d1[159:152];
        7'd21: vec_data_074 = data_d1[167:160];
        7'd22: vec_data_074 = data_d1[175:168];
        7'd23: vec_data_074 = data_d1[183:176];
        7'd24: vec_data_074 = data_d1[191:184];
        7'd25: vec_data_074 = data_d1[199:192];
        7'd26: vec_data_074 = data_d1[207:200];
        7'd27: vec_data_074 = data_d1[215:208];
        7'd28: vec_data_074 = data_d1[223:216];
        7'd29: vec_data_074 = data_d1[231:224];
        7'd30: vec_data_074 = data_d1[239:232];
        7'd31: vec_data_074 = data_d1[247:240];
        7'd32: vec_data_074 = data_d1[255:248];
        7'd33: vec_data_074 = data_d1[263:256];
        7'd34: vec_data_074 = data_d1[271:264];
        7'd35: vec_data_074 = data_d1[279:272];
        7'd36: vec_data_074 = data_d1[287:280];
        7'd37: vec_data_074 = data_d1[295:288];
        7'd38: vec_data_074 = data_d1[303:296];
        7'd39: vec_data_074 = data_d1[311:304];
        7'd40: vec_data_074 = data_d1[319:312];
        7'd41: vec_data_074 = data_d1[327:320];
        7'd42: vec_data_074 = data_d1[335:328];
        7'd43: vec_data_074 = data_d1[343:336];
        7'd44: vec_data_074 = data_d1[351:344];
        7'd45: vec_data_074 = data_d1[359:352];
        7'd46: vec_data_074 = data_d1[367:360];
        7'd47: vec_data_074 = data_d1[375:368];
        7'd48: vec_data_074 = data_d1[383:376];
        7'd49: vec_data_074 = data_d1[391:384];
        7'd50: vec_data_074 = data_d1[399:392];
        7'd51: vec_data_074 = data_d1[407:400];
        7'd52: vec_data_074 = data_d1[415:408];
        7'd53: vec_data_074 = data_d1[423:416];
        7'd54: vec_data_074 = data_d1[431:424];
        7'd55: vec_data_074 = data_d1[439:432];
        7'd56: vec_data_074 = data_d1[447:440];
        7'd57: vec_data_074 = data_d1[455:448];
        7'd58: vec_data_074 = data_d1[463:456];
        7'd59: vec_data_074 = data_d1[471:464];
        7'd60: vec_data_074 = data_d1[479:472];
        7'd61: vec_data_074 = data_d1[487:480];
        7'd62: vec_data_074 = data_d1[495:488];
        7'd63: vec_data_074 = data_d1[503:496];
        7'd64: vec_data_074 = data_d1[511:504];
        7'd65: vec_data_074 = data_d1[519:512];
        7'd66: vec_data_074 = data_d1[527:520];
        7'd67: vec_data_074 = data_d1[535:528];
        7'd68: vec_data_074 = data_d1[543:536];
        7'd69: vec_data_074 = data_d1[551:544];
        7'd70: vec_data_074 = data_d1[559:552];
        7'd71: vec_data_074 = data_d1[567:560];
        7'd72: vec_data_074 = data_d1[575:568];
        7'd73: vec_data_074 = data_d1[583:576];
        7'd74: vec_data_074 = data_d1[591:584];
        7'd75: vec_data_074 = data_d1[599:592];
    endcase
end

always @(
  vec_sum_075_d1
  or data_d1
  ) begin
    vec_data_075 = 8'b0;
    case(vec_sum_075_d1)
        7'd1: vec_data_075 = data_d1[7:0];
        7'd2: vec_data_075 = data_d1[15:8];
        7'd3: vec_data_075 = data_d1[23:16];
        7'd4: vec_data_075 = data_d1[31:24];
        7'd5: vec_data_075 = data_d1[39:32];
        7'd6: vec_data_075 = data_d1[47:40];
        7'd7: vec_data_075 = data_d1[55:48];
        7'd8: vec_data_075 = data_d1[63:56];
        7'd9: vec_data_075 = data_d1[71:64];
        7'd10: vec_data_075 = data_d1[79:72];
        7'd11: vec_data_075 = data_d1[87:80];
        7'd12: vec_data_075 = data_d1[95:88];
        7'd13: vec_data_075 = data_d1[103:96];
        7'd14: vec_data_075 = data_d1[111:104];
        7'd15: vec_data_075 = data_d1[119:112];
        7'd16: vec_data_075 = data_d1[127:120];
        7'd17: vec_data_075 = data_d1[135:128];
        7'd18: vec_data_075 = data_d1[143:136];
        7'd19: vec_data_075 = data_d1[151:144];
        7'd20: vec_data_075 = data_d1[159:152];
        7'd21: vec_data_075 = data_d1[167:160];
        7'd22: vec_data_075 = data_d1[175:168];
        7'd23: vec_data_075 = data_d1[183:176];
        7'd24: vec_data_075 = data_d1[191:184];
        7'd25: vec_data_075 = data_d1[199:192];
        7'd26: vec_data_075 = data_d1[207:200];
        7'd27: vec_data_075 = data_d1[215:208];
        7'd28: vec_data_075 = data_d1[223:216];
        7'd29: vec_data_075 = data_d1[231:224];
        7'd30: vec_data_075 = data_d1[239:232];
        7'd31: vec_data_075 = data_d1[247:240];
        7'd32: vec_data_075 = data_d1[255:248];
        7'd33: vec_data_075 = data_d1[263:256];
        7'd34: vec_data_075 = data_d1[271:264];
        7'd35: vec_data_075 = data_d1[279:272];
        7'd36: vec_data_075 = data_d1[287:280];
        7'd37: vec_data_075 = data_d1[295:288];
        7'd38: vec_data_075 = data_d1[303:296];
        7'd39: vec_data_075 = data_d1[311:304];
        7'd40: vec_data_075 = data_d1[319:312];
        7'd41: vec_data_075 = data_d1[327:320];
        7'd42: vec_data_075 = data_d1[335:328];
        7'd43: vec_data_075 = data_d1[343:336];
        7'd44: vec_data_075 = data_d1[351:344];
        7'd45: vec_data_075 = data_d1[359:352];
        7'd46: vec_data_075 = data_d1[367:360];
        7'd47: vec_data_075 = data_d1[375:368];
        7'd48: vec_data_075 = data_d1[383:376];
        7'd49: vec_data_075 = data_d1[391:384];
        7'd50: vec_data_075 = data_d1[399:392];
        7'd51: vec_data_075 = data_d1[407:400];
        7'd52: vec_data_075 = data_d1[415:408];
        7'd53: vec_data_075 = data_d1[423:416];
        7'd54: vec_data_075 = data_d1[431:424];
        7'd55: vec_data_075 = data_d1[439:432];
        7'd56: vec_data_075 = data_d1[447:440];
        7'd57: vec_data_075 = data_d1[455:448];
        7'd58: vec_data_075 = data_d1[463:456];
        7'd59: vec_data_075 = data_d1[471:464];
        7'd60: vec_data_075 = data_d1[479:472];
        7'd61: vec_data_075 = data_d1[487:480];
        7'd62: vec_data_075 = data_d1[495:488];
        7'd63: vec_data_075 = data_d1[503:496];
        7'd64: vec_data_075 = data_d1[511:504];
        7'd65: vec_data_075 = data_d1[519:512];
        7'd66: vec_data_075 = data_d1[527:520];
        7'd67: vec_data_075 = data_d1[535:528];
        7'd68: vec_data_075 = data_d1[543:536];
        7'd69: vec_data_075 = data_d1[551:544];
        7'd70: vec_data_075 = data_d1[559:552];
        7'd71: vec_data_075 = data_d1[567:560];
        7'd72: vec_data_075 = data_d1[575:568];
        7'd73: vec_data_075 = data_d1[583:576];
        7'd74: vec_data_075 = data_d1[591:584];
        7'd75: vec_data_075 = data_d1[599:592];
        7'd76: vec_data_075 = data_d1[607:600];
    endcase
end

always @(
  vec_sum_076_d1
  or data_d1
  ) begin
    vec_data_076 = 8'b0;
    case(vec_sum_076_d1)
        7'd1: vec_data_076 = data_d1[7:0];
        7'd2: vec_data_076 = data_d1[15:8];
        7'd3: vec_data_076 = data_d1[23:16];
        7'd4: vec_data_076 = data_d1[31:24];
        7'd5: vec_data_076 = data_d1[39:32];
        7'd6: vec_data_076 = data_d1[47:40];
        7'd7: vec_data_076 = data_d1[55:48];
        7'd8: vec_data_076 = data_d1[63:56];
        7'd9: vec_data_076 = data_d1[71:64];
        7'd10: vec_data_076 = data_d1[79:72];
        7'd11: vec_data_076 = data_d1[87:80];
        7'd12: vec_data_076 = data_d1[95:88];
        7'd13: vec_data_076 = data_d1[103:96];
        7'd14: vec_data_076 = data_d1[111:104];
        7'd15: vec_data_076 = data_d1[119:112];
        7'd16: vec_data_076 = data_d1[127:120];
        7'd17: vec_data_076 = data_d1[135:128];
        7'd18: vec_data_076 = data_d1[143:136];
        7'd19: vec_data_076 = data_d1[151:144];
        7'd20: vec_data_076 = data_d1[159:152];
        7'd21: vec_data_076 = data_d1[167:160];
        7'd22: vec_data_076 = data_d1[175:168];
        7'd23: vec_data_076 = data_d1[183:176];
        7'd24: vec_data_076 = data_d1[191:184];
        7'd25: vec_data_076 = data_d1[199:192];
        7'd26: vec_data_076 = data_d1[207:200];
        7'd27: vec_data_076 = data_d1[215:208];
        7'd28: vec_data_076 = data_d1[223:216];
        7'd29: vec_data_076 = data_d1[231:224];
        7'd30: vec_data_076 = data_d1[239:232];
        7'd31: vec_data_076 = data_d1[247:240];
        7'd32: vec_data_076 = data_d1[255:248];
        7'd33: vec_data_076 = data_d1[263:256];
        7'd34: vec_data_076 = data_d1[271:264];
        7'd35: vec_data_076 = data_d1[279:272];
        7'd36: vec_data_076 = data_d1[287:280];
        7'd37: vec_data_076 = data_d1[295:288];
        7'd38: vec_data_076 = data_d1[303:296];
        7'd39: vec_data_076 = data_d1[311:304];
        7'd40: vec_data_076 = data_d1[319:312];
        7'd41: vec_data_076 = data_d1[327:320];
        7'd42: vec_data_076 = data_d1[335:328];
        7'd43: vec_data_076 = data_d1[343:336];
        7'd44: vec_data_076 = data_d1[351:344];
        7'd45: vec_data_076 = data_d1[359:352];
        7'd46: vec_data_076 = data_d1[367:360];
        7'd47: vec_data_076 = data_d1[375:368];
        7'd48: vec_data_076 = data_d1[383:376];
        7'd49: vec_data_076 = data_d1[391:384];
        7'd50: vec_data_076 = data_d1[399:392];
        7'd51: vec_data_076 = data_d1[407:400];
        7'd52: vec_data_076 = data_d1[415:408];
        7'd53: vec_data_076 = data_d1[423:416];
        7'd54: vec_data_076 = data_d1[431:424];
        7'd55: vec_data_076 = data_d1[439:432];
        7'd56: vec_data_076 = data_d1[447:440];
        7'd57: vec_data_076 = data_d1[455:448];
        7'd58: vec_data_076 = data_d1[463:456];
        7'd59: vec_data_076 = data_d1[471:464];
        7'd60: vec_data_076 = data_d1[479:472];
        7'd61: vec_data_076 = data_d1[487:480];
        7'd62: vec_data_076 = data_d1[495:488];
        7'd63: vec_data_076 = data_d1[503:496];
        7'd64: vec_data_076 = data_d1[511:504];
        7'd65: vec_data_076 = data_d1[519:512];
        7'd66: vec_data_076 = data_d1[527:520];
        7'd67: vec_data_076 = data_d1[535:528];
        7'd68: vec_data_076 = data_d1[543:536];
        7'd69: vec_data_076 = data_d1[551:544];
        7'd70: vec_data_076 = data_d1[559:552];
        7'd71: vec_data_076 = data_d1[567:560];
        7'd72: vec_data_076 = data_d1[575:568];
        7'd73: vec_data_076 = data_d1[583:576];
        7'd74: vec_data_076 = data_d1[591:584];
        7'd75: vec_data_076 = data_d1[599:592];
        7'd76: vec_data_076 = data_d1[607:600];
        7'd77: vec_data_076 = data_d1[615:608];
    endcase
end

always @(
  vec_sum_077_d1
  or data_d1
  ) begin
    vec_data_077 = 8'b0;
    case(vec_sum_077_d1)
        7'd1: vec_data_077 = data_d1[7:0];
        7'd2: vec_data_077 = data_d1[15:8];
        7'd3: vec_data_077 = data_d1[23:16];
        7'd4: vec_data_077 = data_d1[31:24];
        7'd5: vec_data_077 = data_d1[39:32];
        7'd6: vec_data_077 = data_d1[47:40];
        7'd7: vec_data_077 = data_d1[55:48];
        7'd8: vec_data_077 = data_d1[63:56];
        7'd9: vec_data_077 = data_d1[71:64];
        7'd10: vec_data_077 = data_d1[79:72];
        7'd11: vec_data_077 = data_d1[87:80];
        7'd12: vec_data_077 = data_d1[95:88];
        7'd13: vec_data_077 = data_d1[103:96];
        7'd14: vec_data_077 = data_d1[111:104];
        7'd15: vec_data_077 = data_d1[119:112];
        7'd16: vec_data_077 = data_d1[127:120];
        7'd17: vec_data_077 = data_d1[135:128];
        7'd18: vec_data_077 = data_d1[143:136];
        7'd19: vec_data_077 = data_d1[151:144];
        7'd20: vec_data_077 = data_d1[159:152];
        7'd21: vec_data_077 = data_d1[167:160];
        7'd22: vec_data_077 = data_d1[175:168];
        7'd23: vec_data_077 = data_d1[183:176];
        7'd24: vec_data_077 = data_d1[191:184];
        7'd25: vec_data_077 = data_d1[199:192];
        7'd26: vec_data_077 = data_d1[207:200];
        7'd27: vec_data_077 = data_d1[215:208];
        7'd28: vec_data_077 = data_d1[223:216];
        7'd29: vec_data_077 = data_d1[231:224];
        7'd30: vec_data_077 = data_d1[239:232];
        7'd31: vec_data_077 = data_d1[247:240];
        7'd32: vec_data_077 = data_d1[255:248];
        7'd33: vec_data_077 = data_d1[263:256];
        7'd34: vec_data_077 = data_d1[271:264];
        7'd35: vec_data_077 = data_d1[279:272];
        7'd36: vec_data_077 = data_d1[287:280];
        7'd37: vec_data_077 = data_d1[295:288];
        7'd38: vec_data_077 = data_d1[303:296];
        7'd39: vec_data_077 = data_d1[311:304];
        7'd40: vec_data_077 = data_d1[319:312];
        7'd41: vec_data_077 = data_d1[327:320];
        7'd42: vec_data_077 = data_d1[335:328];
        7'd43: vec_data_077 = data_d1[343:336];
        7'd44: vec_data_077 = data_d1[351:344];
        7'd45: vec_data_077 = data_d1[359:352];
        7'd46: vec_data_077 = data_d1[367:360];
        7'd47: vec_data_077 = data_d1[375:368];
        7'd48: vec_data_077 = data_d1[383:376];
        7'd49: vec_data_077 = data_d1[391:384];
        7'd50: vec_data_077 = data_d1[399:392];
        7'd51: vec_data_077 = data_d1[407:400];
        7'd52: vec_data_077 = data_d1[415:408];
        7'd53: vec_data_077 = data_d1[423:416];
        7'd54: vec_data_077 = data_d1[431:424];
        7'd55: vec_data_077 = data_d1[439:432];
        7'd56: vec_data_077 = data_d1[447:440];
        7'd57: vec_data_077 = data_d1[455:448];
        7'd58: vec_data_077 = data_d1[463:456];
        7'd59: vec_data_077 = data_d1[471:464];
        7'd60: vec_data_077 = data_d1[479:472];
        7'd61: vec_data_077 = data_d1[487:480];
        7'd62: vec_data_077 = data_d1[495:488];
        7'd63: vec_data_077 = data_d1[503:496];
        7'd64: vec_data_077 = data_d1[511:504];
        7'd65: vec_data_077 = data_d1[519:512];
        7'd66: vec_data_077 = data_d1[527:520];
        7'd67: vec_data_077 = data_d1[535:528];
        7'd68: vec_data_077 = data_d1[543:536];
        7'd69: vec_data_077 = data_d1[551:544];
        7'd70: vec_data_077 = data_d1[559:552];
        7'd71: vec_data_077 = data_d1[567:560];
        7'd72: vec_data_077 = data_d1[575:568];
        7'd73: vec_data_077 = data_d1[583:576];
        7'd74: vec_data_077 = data_d1[591:584];
        7'd75: vec_data_077 = data_d1[599:592];
        7'd76: vec_data_077 = data_d1[607:600];
        7'd77: vec_data_077 = data_d1[615:608];
        7'd78: vec_data_077 = data_d1[623:616];
    endcase
end

always @(
  vec_sum_078_d1
  or data_d1
  ) begin
    vec_data_078 = 8'b0;
    case(vec_sum_078_d1)
        7'd1: vec_data_078 = data_d1[7:0];
        7'd2: vec_data_078 = data_d1[15:8];
        7'd3: vec_data_078 = data_d1[23:16];
        7'd4: vec_data_078 = data_d1[31:24];
        7'd5: vec_data_078 = data_d1[39:32];
        7'd6: vec_data_078 = data_d1[47:40];
        7'd7: vec_data_078 = data_d1[55:48];
        7'd8: vec_data_078 = data_d1[63:56];
        7'd9: vec_data_078 = data_d1[71:64];
        7'd10: vec_data_078 = data_d1[79:72];
        7'd11: vec_data_078 = data_d1[87:80];
        7'd12: vec_data_078 = data_d1[95:88];
        7'd13: vec_data_078 = data_d1[103:96];
        7'd14: vec_data_078 = data_d1[111:104];
        7'd15: vec_data_078 = data_d1[119:112];
        7'd16: vec_data_078 = data_d1[127:120];
        7'd17: vec_data_078 = data_d1[135:128];
        7'd18: vec_data_078 = data_d1[143:136];
        7'd19: vec_data_078 = data_d1[151:144];
        7'd20: vec_data_078 = data_d1[159:152];
        7'd21: vec_data_078 = data_d1[167:160];
        7'd22: vec_data_078 = data_d1[175:168];
        7'd23: vec_data_078 = data_d1[183:176];
        7'd24: vec_data_078 = data_d1[191:184];
        7'd25: vec_data_078 = data_d1[199:192];
        7'd26: vec_data_078 = data_d1[207:200];
        7'd27: vec_data_078 = data_d1[215:208];
        7'd28: vec_data_078 = data_d1[223:216];
        7'd29: vec_data_078 = data_d1[231:224];
        7'd30: vec_data_078 = data_d1[239:232];
        7'd31: vec_data_078 = data_d1[247:240];
        7'd32: vec_data_078 = data_d1[255:248];
        7'd33: vec_data_078 = data_d1[263:256];
        7'd34: vec_data_078 = data_d1[271:264];
        7'd35: vec_data_078 = data_d1[279:272];
        7'd36: vec_data_078 = data_d1[287:280];
        7'd37: vec_data_078 = data_d1[295:288];
        7'd38: vec_data_078 = data_d1[303:296];
        7'd39: vec_data_078 = data_d1[311:304];
        7'd40: vec_data_078 = data_d1[319:312];
        7'd41: vec_data_078 = data_d1[327:320];
        7'd42: vec_data_078 = data_d1[335:328];
        7'd43: vec_data_078 = data_d1[343:336];
        7'd44: vec_data_078 = data_d1[351:344];
        7'd45: vec_data_078 = data_d1[359:352];
        7'd46: vec_data_078 = data_d1[367:360];
        7'd47: vec_data_078 = data_d1[375:368];
        7'd48: vec_data_078 = data_d1[383:376];
        7'd49: vec_data_078 = data_d1[391:384];
        7'd50: vec_data_078 = data_d1[399:392];
        7'd51: vec_data_078 = data_d1[407:400];
        7'd52: vec_data_078 = data_d1[415:408];
        7'd53: vec_data_078 = data_d1[423:416];
        7'd54: vec_data_078 = data_d1[431:424];
        7'd55: vec_data_078 = data_d1[439:432];
        7'd56: vec_data_078 = data_d1[447:440];
        7'd57: vec_data_078 = data_d1[455:448];
        7'd58: vec_data_078 = data_d1[463:456];
        7'd59: vec_data_078 = data_d1[471:464];
        7'd60: vec_data_078 = data_d1[479:472];
        7'd61: vec_data_078 = data_d1[487:480];
        7'd62: vec_data_078 = data_d1[495:488];
        7'd63: vec_data_078 = data_d1[503:496];
        7'd64: vec_data_078 = data_d1[511:504];
        7'd65: vec_data_078 = data_d1[519:512];
        7'd66: vec_data_078 = data_d1[527:520];
        7'd67: vec_data_078 = data_d1[535:528];
        7'd68: vec_data_078 = data_d1[543:536];
        7'd69: vec_data_078 = data_d1[551:544];
        7'd70: vec_data_078 = data_d1[559:552];
        7'd71: vec_data_078 = data_d1[567:560];
        7'd72: vec_data_078 = data_d1[575:568];
        7'd73: vec_data_078 = data_d1[583:576];
        7'd74: vec_data_078 = data_d1[591:584];
        7'd75: vec_data_078 = data_d1[599:592];
        7'd76: vec_data_078 = data_d1[607:600];
        7'd77: vec_data_078 = data_d1[615:608];
        7'd78: vec_data_078 = data_d1[623:616];
        7'd79: vec_data_078 = data_d1[631:624];
    endcase
end

always @(
  vec_sum_079_d1
  or data_d1
  ) begin
    vec_data_079 = 8'b0;
    case(vec_sum_079_d1)
        7'd1: vec_data_079 = data_d1[7:0];
        7'd2: vec_data_079 = data_d1[15:8];
        7'd3: vec_data_079 = data_d1[23:16];
        7'd4: vec_data_079 = data_d1[31:24];
        7'd5: vec_data_079 = data_d1[39:32];
        7'd6: vec_data_079 = data_d1[47:40];
        7'd7: vec_data_079 = data_d1[55:48];
        7'd8: vec_data_079 = data_d1[63:56];
        7'd9: vec_data_079 = data_d1[71:64];
        7'd10: vec_data_079 = data_d1[79:72];
        7'd11: vec_data_079 = data_d1[87:80];
        7'd12: vec_data_079 = data_d1[95:88];
        7'd13: vec_data_079 = data_d1[103:96];
        7'd14: vec_data_079 = data_d1[111:104];
        7'd15: vec_data_079 = data_d1[119:112];
        7'd16: vec_data_079 = data_d1[127:120];
        7'd17: vec_data_079 = data_d1[135:128];
        7'd18: vec_data_079 = data_d1[143:136];
        7'd19: vec_data_079 = data_d1[151:144];
        7'd20: vec_data_079 = data_d1[159:152];
        7'd21: vec_data_079 = data_d1[167:160];
        7'd22: vec_data_079 = data_d1[175:168];
        7'd23: vec_data_079 = data_d1[183:176];
        7'd24: vec_data_079 = data_d1[191:184];
        7'd25: vec_data_079 = data_d1[199:192];
        7'd26: vec_data_079 = data_d1[207:200];
        7'd27: vec_data_079 = data_d1[215:208];
        7'd28: vec_data_079 = data_d1[223:216];
        7'd29: vec_data_079 = data_d1[231:224];
        7'd30: vec_data_079 = data_d1[239:232];
        7'd31: vec_data_079 = data_d1[247:240];
        7'd32: vec_data_079 = data_d1[255:248];
        7'd33: vec_data_079 = data_d1[263:256];
        7'd34: vec_data_079 = data_d1[271:264];
        7'd35: vec_data_079 = data_d1[279:272];
        7'd36: vec_data_079 = data_d1[287:280];
        7'd37: vec_data_079 = data_d1[295:288];
        7'd38: vec_data_079 = data_d1[303:296];
        7'd39: vec_data_079 = data_d1[311:304];
        7'd40: vec_data_079 = data_d1[319:312];
        7'd41: vec_data_079 = data_d1[327:320];
        7'd42: vec_data_079 = data_d1[335:328];
        7'd43: vec_data_079 = data_d1[343:336];
        7'd44: vec_data_079 = data_d1[351:344];
        7'd45: vec_data_079 = data_d1[359:352];
        7'd46: vec_data_079 = data_d1[367:360];
        7'd47: vec_data_079 = data_d1[375:368];
        7'd48: vec_data_079 = data_d1[383:376];
        7'd49: vec_data_079 = data_d1[391:384];
        7'd50: vec_data_079 = data_d1[399:392];
        7'd51: vec_data_079 = data_d1[407:400];
        7'd52: vec_data_079 = data_d1[415:408];
        7'd53: vec_data_079 = data_d1[423:416];
        7'd54: vec_data_079 = data_d1[431:424];
        7'd55: vec_data_079 = data_d1[439:432];
        7'd56: vec_data_079 = data_d1[447:440];
        7'd57: vec_data_079 = data_d1[455:448];
        7'd58: vec_data_079 = data_d1[463:456];
        7'd59: vec_data_079 = data_d1[471:464];
        7'd60: vec_data_079 = data_d1[479:472];
        7'd61: vec_data_079 = data_d1[487:480];
        7'd62: vec_data_079 = data_d1[495:488];
        7'd63: vec_data_079 = data_d1[503:496];
        7'd64: vec_data_079 = data_d1[511:504];
        7'd65: vec_data_079 = data_d1[519:512];
        7'd66: vec_data_079 = data_d1[527:520];
        7'd67: vec_data_079 = data_d1[535:528];
        7'd68: vec_data_079 = data_d1[543:536];
        7'd69: vec_data_079 = data_d1[551:544];
        7'd70: vec_data_079 = data_d1[559:552];
        7'd71: vec_data_079 = data_d1[567:560];
        7'd72: vec_data_079 = data_d1[575:568];
        7'd73: vec_data_079 = data_d1[583:576];
        7'd74: vec_data_079 = data_d1[591:584];
        7'd75: vec_data_079 = data_d1[599:592];
        7'd76: vec_data_079 = data_d1[607:600];
        7'd77: vec_data_079 = data_d1[615:608];
        7'd78: vec_data_079 = data_d1[623:616];
        7'd79: vec_data_079 = data_d1[631:624];
        7'd80: vec_data_079 = data_d1[639:632];
    endcase
end

always @(
  vec_sum_080_d1
  or data_d1
  ) begin
    vec_data_080 = 8'b0;
    case(vec_sum_080_d1)
        7'd1: vec_data_080 = data_d1[7:0];
        7'd2: vec_data_080 = data_d1[15:8];
        7'd3: vec_data_080 = data_d1[23:16];
        7'd4: vec_data_080 = data_d1[31:24];
        7'd5: vec_data_080 = data_d1[39:32];
        7'd6: vec_data_080 = data_d1[47:40];
        7'd7: vec_data_080 = data_d1[55:48];
        7'd8: vec_data_080 = data_d1[63:56];
        7'd9: vec_data_080 = data_d1[71:64];
        7'd10: vec_data_080 = data_d1[79:72];
        7'd11: vec_data_080 = data_d1[87:80];
        7'd12: vec_data_080 = data_d1[95:88];
        7'd13: vec_data_080 = data_d1[103:96];
        7'd14: vec_data_080 = data_d1[111:104];
        7'd15: vec_data_080 = data_d1[119:112];
        7'd16: vec_data_080 = data_d1[127:120];
        7'd17: vec_data_080 = data_d1[135:128];
        7'd18: vec_data_080 = data_d1[143:136];
        7'd19: vec_data_080 = data_d1[151:144];
        7'd20: vec_data_080 = data_d1[159:152];
        7'd21: vec_data_080 = data_d1[167:160];
        7'd22: vec_data_080 = data_d1[175:168];
        7'd23: vec_data_080 = data_d1[183:176];
        7'd24: vec_data_080 = data_d1[191:184];
        7'd25: vec_data_080 = data_d1[199:192];
        7'd26: vec_data_080 = data_d1[207:200];
        7'd27: vec_data_080 = data_d1[215:208];
        7'd28: vec_data_080 = data_d1[223:216];
        7'd29: vec_data_080 = data_d1[231:224];
        7'd30: vec_data_080 = data_d1[239:232];
        7'd31: vec_data_080 = data_d1[247:240];
        7'd32: vec_data_080 = data_d1[255:248];
        7'd33: vec_data_080 = data_d1[263:256];
        7'd34: vec_data_080 = data_d1[271:264];
        7'd35: vec_data_080 = data_d1[279:272];
        7'd36: vec_data_080 = data_d1[287:280];
        7'd37: vec_data_080 = data_d1[295:288];
        7'd38: vec_data_080 = data_d1[303:296];
        7'd39: vec_data_080 = data_d1[311:304];
        7'd40: vec_data_080 = data_d1[319:312];
        7'd41: vec_data_080 = data_d1[327:320];
        7'd42: vec_data_080 = data_d1[335:328];
        7'd43: vec_data_080 = data_d1[343:336];
        7'd44: vec_data_080 = data_d1[351:344];
        7'd45: vec_data_080 = data_d1[359:352];
        7'd46: vec_data_080 = data_d1[367:360];
        7'd47: vec_data_080 = data_d1[375:368];
        7'd48: vec_data_080 = data_d1[383:376];
        7'd49: vec_data_080 = data_d1[391:384];
        7'd50: vec_data_080 = data_d1[399:392];
        7'd51: vec_data_080 = data_d1[407:400];
        7'd52: vec_data_080 = data_d1[415:408];
        7'd53: vec_data_080 = data_d1[423:416];
        7'd54: vec_data_080 = data_d1[431:424];
        7'd55: vec_data_080 = data_d1[439:432];
        7'd56: vec_data_080 = data_d1[447:440];
        7'd57: vec_data_080 = data_d1[455:448];
        7'd58: vec_data_080 = data_d1[463:456];
        7'd59: vec_data_080 = data_d1[471:464];
        7'd60: vec_data_080 = data_d1[479:472];
        7'd61: vec_data_080 = data_d1[487:480];
        7'd62: vec_data_080 = data_d1[495:488];
        7'd63: vec_data_080 = data_d1[503:496];
        7'd64: vec_data_080 = data_d1[511:504];
        7'd65: vec_data_080 = data_d1[519:512];
        7'd66: vec_data_080 = data_d1[527:520];
        7'd67: vec_data_080 = data_d1[535:528];
        7'd68: vec_data_080 = data_d1[543:536];
        7'd69: vec_data_080 = data_d1[551:544];
        7'd70: vec_data_080 = data_d1[559:552];
        7'd71: vec_data_080 = data_d1[567:560];
        7'd72: vec_data_080 = data_d1[575:568];
        7'd73: vec_data_080 = data_d1[583:576];
        7'd74: vec_data_080 = data_d1[591:584];
        7'd75: vec_data_080 = data_d1[599:592];
        7'd76: vec_data_080 = data_d1[607:600];
        7'd77: vec_data_080 = data_d1[615:608];
        7'd78: vec_data_080 = data_d1[623:616];
        7'd79: vec_data_080 = data_d1[631:624];
        7'd80: vec_data_080 = data_d1[639:632];
        7'd81: vec_data_080 = data_d1[647:640];
    endcase
end

always @(
  vec_sum_081_d1
  or data_d1
  ) begin
    vec_data_081 = 8'b0;
    case(vec_sum_081_d1)
        7'd1: vec_data_081 = data_d1[7:0];
        7'd2: vec_data_081 = data_d1[15:8];
        7'd3: vec_data_081 = data_d1[23:16];
        7'd4: vec_data_081 = data_d1[31:24];
        7'd5: vec_data_081 = data_d1[39:32];
        7'd6: vec_data_081 = data_d1[47:40];
        7'd7: vec_data_081 = data_d1[55:48];
        7'd8: vec_data_081 = data_d1[63:56];
        7'd9: vec_data_081 = data_d1[71:64];
        7'd10: vec_data_081 = data_d1[79:72];
        7'd11: vec_data_081 = data_d1[87:80];
        7'd12: vec_data_081 = data_d1[95:88];
        7'd13: vec_data_081 = data_d1[103:96];
        7'd14: vec_data_081 = data_d1[111:104];
        7'd15: vec_data_081 = data_d1[119:112];
        7'd16: vec_data_081 = data_d1[127:120];
        7'd17: vec_data_081 = data_d1[135:128];
        7'd18: vec_data_081 = data_d1[143:136];
        7'd19: vec_data_081 = data_d1[151:144];
        7'd20: vec_data_081 = data_d1[159:152];
        7'd21: vec_data_081 = data_d1[167:160];
        7'd22: vec_data_081 = data_d1[175:168];
        7'd23: vec_data_081 = data_d1[183:176];
        7'd24: vec_data_081 = data_d1[191:184];
        7'd25: vec_data_081 = data_d1[199:192];
        7'd26: vec_data_081 = data_d1[207:200];
        7'd27: vec_data_081 = data_d1[215:208];
        7'd28: vec_data_081 = data_d1[223:216];
        7'd29: vec_data_081 = data_d1[231:224];
        7'd30: vec_data_081 = data_d1[239:232];
        7'd31: vec_data_081 = data_d1[247:240];
        7'd32: vec_data_081 = data_d1[255:248];
        7'd33: vec_data_081 = data_d1[263:256];
        7'd34: vec_data_081 = data_d1[271:264];
        7'd35: vec_data_081 = data_d1[279:272];
        7'd36: vec_data_081 = data_d1[287:280];
        7'd37: vec_data_081 = data_d1[295:288];
        7'd38: vec_data_081 = data_d1[303:296];
        7'd39: vec_data_081 = data_d1[311:304];
        7'd40: vec_data_081 = data_d1[319:312];
        7'd41: vec_data_081 = data_d1[327:320];
        7'd42: vec_data_081 = data_d1[335:328];
        7'd43: vec_data_081 = data_d1[343:336];
        7'd44: vec_data_081 = data_d1[351:344];
        7'd45: vec_data_081 = data_d1[359:352];
        7'd46: vec_data_081 = data_d1[367:360];
        7'd47: vec_data_081 = data_d1[375:368];
        7'd48: vec_data_081 = data_d1[383:376];
        7'd49: vec_data_081 = data_d1[391:384];
        7'd50: vec_data_081 = data_d1[399:392];
        7'd51: vec_data_081 = data_d1[407:400];
        7'd52: vec_data_081 = data_d1[415:408];
        7'd53: vec_data_081 = data_d1[423:416];
        7'd54: vec_data_081 = data_d1[431:424];
        7'd55: vec_data_081 = data_d1[439:432];
        7'd56: vec_data_081 = data_d1[447:440];
        7'd57: vec_data_081 = data_d1[455:448];
        7'd58: vec_data_081 = data_d1[463:456];
        7'd59: vec_data_081 = data_d1[471:464];
        7'd60: vec_data_081 = data_d1[479:472];
        7'd61: vec_data_081 = data_d1[487:480];
        7'd62: vec_data_081 = data_d1[495:488];
        7'd63: vec_data_081 = data_d1[503:496];
        7'd64: vec_data_081 = data_d1[511:504];
        7'd65: vec_data_081 = data_d1[519:512];
        7'd66: vec_data_081 = data_d1[527:520];
        7'd67: vec_data_081 = data_d1[535:528];
        7'd68: vec_data_081 = data_d1[543:536];
        7'd69: vec_data_081 = data_d1[551:544];
        7'd70: vec_data_081 = data_d1[559:552];
        7'd71: vec_data_081 = data_d1[567:560];
        7'd72: vec_data_081 = data_d1[575:568];
        7'd73: vec_data_081 = data_d1[583:576];
        7'd74: vec_data_081 = data_d1[591:584];
        7'd75: vec_data_081 = data_d1[599:592];
        7'd76: vec_data_081 = data_d1[607:600];
        7'd77: vec_data_081 = data_d1[615:608];
        7'd78: vec_data_081 = data_d1[623:616];
        7'd79: vec_data_081 = data_d1[631:624];
        7'd80: vec_data_081 = data_d1[639:632];
        7'd81: vec_data_081 = data_d1[647:640];
        7'd82: vec_data_081 = data_d1[655:648];
    endcase
end

always @(
  vec_sum_082_d1
  or data_d1
  ) begin
    vec_data_082 = 8'b0;
    case(vec_sum_082_d1)
        7'd1: vec_data_082 = data_d1[7:0];
        7'd2: vec_data_082 = data_d1[15:8];
        7'd3: vec_data_082 = data_d1[23:16];
        7'd4: vec_data_082 = data_d1[31:24];
        7'd5: vec_data_082 = data_d1[39:32];
        7'd6: vec_data_082 = data_d1[47:40];
        7'd7: vec_data_082 = data_d1[55:48];
        7'd8: vec_data_082 = data_d1[63:56];
        7'd9: vec_data_082 = data_d1[71:64];
        7'd10: vec_data_082 = data_d1[79:72];
        7'd11: vec_data_082 = data_d1[87:80];
        7'd12: vec_data_082 = data_d1[95:88];
        7'd13: vec_data_082 = data_d1[103:96];
        7'd14: vec_data_082 = data_d1[111:104];
        7'd15: vec_data_082 = data_d1[119:112];
        7'd16: vec_data_082 = data_d1[127:120];
        7'd17: vec_data_082 = data_d1[135:128];
        7'd18: vec_data_082 = data_d1[143:136];
        7'd19: vec_data_082 = data_d1[151:144];
        7'd20: vec_data_082 = data_d1[159:152];
        7'd21: vec_data_082 = data_d1[167:160];
        7'd22: vec_data_082 = data_d1[175:168];
        7'd23: vec_data_082 = data_d1[183:176];
        7'd24: vec_data_082 = data_d1[191:184];
        7'd25: vec_data_082 = data_d1[199:192];
        7'd26: vec_data_082 = data_d1[207:200];
        7'd27: vec_data_082 = data_d1[215:208];
        7'd28: vec_data_082 = data_d1[223:216];
        7'd29: vec_data_082 = data_d1[231:224];
        7'd30: vec_data_082 = data_d1[239:232];
        7'd31: vec_data_082 = data_d1[247:240];
        7'd32: vec_data_082 = data_d1[255:248];
        7'd33: vec_data_082 = data_d1[263:256];
        7'd34: vec_data_082 = data_d1[271:264];
        7'd35: vec_data_082 = data_d1[279:272];
        7'd36: vec_data_082 = data_d1[287:280];
        7'd37: vec_data_082 = data_d1[295:288];
        7'd38: vec_data_082 = data_d1[303:296];
        7'd39: vec_data_082 = data_d1[311:304];
        7'd40: vec_data_082 = data_d1[319:312];
        7'd41: vec_data_082 = data_d1[327:320];
        7'd42: vec_data_082 = data_d1[335:328];
        7'd43: vec_data_082 = data_d1[343:336];
        7'd44: vec_data_082 = data_d1[351:344];
        7'd45: vec_data_082 = data_d1[359:352];
        7'd46: vec_data_082 = data_d1[367:360];
        7'd47: vec_data_082 = data_d1[375:368];
        7'd48: vec_data_082 = data_d1[383:376];
        7'd49: vec_data_082 = data_d1[391:384];
        7'd50: vec_data_082 = data_d1[399:392];
        7'd51: vec_data_082 = data_d1[407:400];
        7'd52: vec_data_082 = data_d1[415:408];
        7'd53: vec_data_082 = data_d1[423:416];
        7'd54: vec_data_082 = data_d1[431:424];
        7'd55: vec_data_082 = data_d1[439:432];
        7'd56: vec_data_082 = data_d1[447:440];
        7'd57: vec_data_082 = data_d1[455:448];
        7'd58: vec_data_082 = data_d1[463:456];
        7'd59: vec_data_082 = data_d1[471:464];
        7'd60: vec_data_082 = data_d1[479:472];
        7'd61: vec_data_082 = data_d1[487:480];
        7'd62: vec_data_082 = data_d1[495:488];
        7'd63: vec_data_082 = data_d1[503:496];
        7'd64: vec_data_082 = data_d1[511:504];
        7'd65: vec_data_082 = data_d1[519:512];
        7'd66: vec_data_082 = data_d1[527:520];
        7'd67: vec_data_082 = data_d1[535:528];
        7'd68: vec_data_082 = data_d1[543:536];
        7'd69: vec_data_082 = data_d1[551:544];
        7'd70: vec_data_082 = data_d1[559:552];
        7'd71: vec_data_082 = data_d1[567:560];
        7'd72: vec_data_082 = data_d1[575:568];
        7'd73: vec_data_082 = data_d1[583:576];
        7'd74: vec_data_082 = data_d1[591:584];
        7'd75: vec_data_082 = data_d1[599:592];
        7'd76: vec_data_082 = data_d1[607:600];
        7'd77: vec_data_082 = data_d1[615:608];
        7'd78: vec_data_082 = data_d1[623:616];
        7'd79: vec_data_082 = data_d1[631:624];
        7'd80: vec_data_082 = data_d1[639:632];
        7'd81: vec_data_082 = data_d1[647:640];
        7'd82: vec_data_082 = data_d1[655:648];
        7'd83: vec_data_082 = data_d1[663:656];
    endcase
end

always @(
  vec_sum_083_d1
  or data_d1
  ) begin
    vec_data_083 = 8'b0;
    case(vec_sum_083_d1)
        7'd1: vec_data_083 = data_d1[7:0];
        7'd2: vec_data_083 = data_d1[15:8];
        7'd3: vec_data_083 = data_d1[23:16];
        7'd4: vec_data_083 = data_d1[31:24];
        7'd5: vec_data_083 = data_d1[39:32];
        7'd6: vec_data_083 = data_d1[47:40];
        7'd7: vec_data_083 = data_d1[55:48];
        7'd8: vec_data_083 = data_d1[63:56];
        7'd9: vec_data_083 = data_d1[71:64];
        7'd10: vec_data_083 = data_d1[79:72];
        7'd11: vec_data_083 = data_d1[87:80];
        7'd12: vec_data_083 = data_d1[95:88];
        7'd13: vec_data_083 = data_d1[103:96];
        7'd14: vec_data_083 = data_d1[111:104];
        7'd15: vec_data_083 = data_d1[119:112];
        7'd16: vec_data_083 = data_d1[127:120];
        7'd17: vec_data_083 = data_d1[135:128];
        7'd18: vec_data_083 = data_d1[143:136];
        7'd19: vec_data_083 = data_d1[151:144];
        7'd20: vec_data_083 = data_d1[159:152];
        7'd21: vec_data_083 = data_d1[167:160];
        7'd22: vec_data_083 = data_d1[175:168];
        7'd23: vec_data_083 = data_d1[183:176];
        7'd24: vec_data_083 = data_d1[191:184];
        7'd25: vec_data_083 = data_d1[199:192];
        7'd26: vec_data_083 = data_d1[207:200];
        7'd27: vec_data_083 = data_d1[215:208];
        7'd28: vec_data_083 = data_d1[223:216];
        7'd29: vec_data_083 = data_d1[231:224];
        7'd30: vec_data_083 = data_d1[239:232];
        7'd31: vec_data_083 = data_d1[247:240];
        7'd32: vec_data_083 = data_d1[255:248];
        7'd33: vec_data_083 = data_d1[263:256];
        7'd34: vec_data_083 = data_d1[271:264];
        7'd35: vec_data_083 = data_d1[279:272];
        7'd36: vec_data_083 = data_d1[287:280];
        7'd37: vec_data_083 = data_d1[295:288];
        7'd38: vec_data_083 = data_d1[303:296];
        7'd39: vec_data_083 = data_d1[311:304];
        7'd40: vec_data_083 = data_d1[319:312];
        7'd41: vec_data_083 = data_d1[327:320];
        7'd42: vec_data_083 = data_d1[335:328];
        7'd43: vec_data_083 = data_d1[343:336];
        7'd44: vec_data_083 = data_d1[351:344];
        7'd45: vec_data_083 = data_d1[359:352];
        7'd46: vec_data_083 = data_d1[367:360];
        7'd47: vec_data_083 = data_d1[375:368];
        7'd48: vec_data_083 = data_d1[383:376];
        7'd49: vec_data_083 = data_d1[391:384];
        7'd50: vec_data_083 = data_d1[399:392];
        7'd51: vec_data_083 = data_d1[407:400];
        7'd52: vec_data_083 = data_d1[415:408];
        7'd53: vec_data_083 = data_d1[423:416];
        7'd54: vec_data_083 = data_d1[431:424];
        7'd55: vec_data_083 = data_d1[439:432];
        7'd56: vec_data_083 = data_d1[447:440];
        7'd57: vec_data_083 = data_d1[455:448];
        7'd58: vec_data_083 = data_d1[463:456];
        7'd59: vec_data_083 = data_d1[471:464];
        7'd60: vec_data_083 = data_d1[479:472];
        7'd61: vec_data_083 = data_d1[487:480];
        7'd62: vec_data_083 = data_d1[495:488];
        7'd63: vec_data_083 = data_d1[503:496];
        7'd64: vec_data_083 = data_d1[511:504];
        7'd65: vec_data_083 = data_d1[519:512];
        7'd66: vec_data_083 = data_d1[527:520];
        7'd67: vec_data_083 = data_d1[535:528];
        7'd68: vec_data_083 = data_d1[543:536];
        7'd69: vec_data_083 = data_d1[551:544];
        7'd70: vec_data_083 = data_d1[559:552];
        7'd71: vec_data_083 = data_d1[567:560];
        7'd72: vec_data_083 = data_d1[575:568];
        7'd73: vec_data_083 = data_d1[583:576];
        7'd74: vec_data_083 = data_d1[591:584];
        7'd75: vec_data_083 = data_d1[599:592];
        7'd76: vec_data_083 = data_d1[607:600];
        7'd77: vec_data_083 = data_d1[615:608];
        7'd78: vec_data_083 = data_d1[623:616];
        7'd79: vec_data_083 = data_d1[631:624];
        7'd80: vec_data_083 = data_d1[639:632];
        7'd81: vec_data_083 = data_d1[647:640];
        7'd82: vec_data_083 = data_d1[655:648];
        7'd83: vec_data_083 = data_d1[663:656];
        7'd84: vec_data_083 = data_d1[671:664];
    endcase
end

always @(
  vec_sum_084_d1
  or data_d1
  ) begin
    vec_data_084 = 8'b0;
    case(vec_sum_084_d1)
        7'd1: vec_data_084 = data_d1[7:0];
        7'd2: vec_data_084 = data_d1[15:8];
        7'd3: vec_data_084 = data_d1[23:16];
        7'd4: vec_data_084 = data_d1[31:24];
        7'd5: vec_data_084 = data_d1[39:32];
        7'd6: vec_data_084 = data_d1[47:40];
        7'd7: vec_data_084 = data_d1[55:48];
        7'd8: vec_data_084 = data_d1[63:56];
        7'd9: vec_data_084 = data_d1[71:64];
        7'd10: vec_data_084 = data_d1[79:72];
        7'd11: vec_data_084 = data_d1[87:80];
        7'd12: vec_data_084 = data_d1[95:88];
        7'd13: vec_data_084 = data_d1[103:96];
        7'd14: vec_data_084 = data_d1[111:104];
        7'd15: vec_data_084 = data_d1[119:112];
        7'd16: vec_data_084 = data_d1[127:120];
        7'd17: vec_data_084 = data_d1[135:128];
        7'd18: vec_data_084 = data_d1[143:136];
        7'd19: vec_data_084 = data_d1[151:144];
        7'd20: vec_data_084 = data_d1[159:152];
        7'd21: vec_data_084 = data_d1[167:160];
        7'd22: vec_data_084 = data_d1[175:168];
        7'd23: vec_data_084 = data_d1[183:176];
        7'd24: vec_data_084 = data_d1[191:184];
        7'd25: vec_data_084 = data_d1[199:192];
        7'd26: vec_data_084 = data_d1[207:200];
        7'd27: vec_data_084 = data_d1[215:208];
        7'd28: vec_data_084 = data_d1[223:216];
        7'd29: vec_data_084 = data_d1[231:224];
        7'd30: vec_data_084 = data_d1[239:232];
        7'd31: vec_data_084 = data_d1[247:240];
        7'd32: vec_data_084 = data_d1[255:248];
        7'd33: vec_data_084 = data_d1[263:256];
        7'd34: vec_data_084 = data_d1[271:264];
        7'd35: vec_data_084 = data_d1[279:272];
        7'd36: vec_data_084 = data_d1[287:280];
        7'd37: vec_data_084 = data_d1[295:288];
        7'd38: vec_data_084 = data_d1[303:296];
        7'd39: vec_data_084 = data_d1[311:304];
        7'd40: vec_data_084 = data_d1[319:312];
        7'd41: vec_data_084 = data_d1[327:320];
        7'd42: vec_data_084 = data_d1[335:328];
        7'd43: vec_data_084 = data_d1[343:336];
        7'd44: vec_data_084 = data_d1[351:344];
        7'd45: vec_data_084 = data_d1[359:352];
        7'd46: vec_data_084 = data_d1[367:360];
        7'd47: vec_data_084 = data_d1[375:368];
        7'd48: vec_data_084 = data_d1[383:376];
        7'd49: vec_data_084 = data_d1[391:384];
        7'd50: vec_data_084 = data_d1[399:392];
        7'd51: vec_data_084 = data_d1[407:400];
        7'd52: vec_data_084 = data_d1[415:408];
        7'd53: vec_data_084 = data_d1[423:416];
        7'd54: vec_data_084 = data_d1[431:424];
        7'd55: vec_data_084 = data_d1[439:432];
        7'd56: vec_data_084 = data_d1[447:440];
        7'd57: vec_data_084 = data_d1[455:448];
        7'd58: vec_data_084 = data_d1[463:456];
        7'd59: vec_data_084 = data_d1[471:464];
        7'd60: vec_data_084 = data_d1[479:472];
        7'd61: vec_data_084 = data_d1[487:480];
        7'd62: vec_data_084 = data_d1[495:488];
        7'd63: vec_data_084 = data_d1[503:496];
        7'd64: vec_data_084 = data_d1[511:504];
        7'd65: vec_data_084 = data_d1[519:512];
        7'd66: vec_data_084 = data_d1[527:520];
        7'd67: vec_data_084 = data_d1[535:528];
        7'd68: vec_data_084 = data_d1[543:536];
        7'd69: vec_data_084 = data_d1[551:544];
        7'd70: vec_data_084 = data_d1[559:552];
        7'd71: vec_data_084 = data_d1[567:560];
        7'd72: vec_data_084 = data_d1[575:568];
        7'd73: vec_data_084 = data_d1[583:576];
        7'd74: vec_data_084 = data_d1[591:584];
        7'd75: vec_data_084 = data_d1[599:592];
        7'd76: vec_data_084 = data_d1[607:600];
        7'd77: vec_data_084 = data_d1[615:608];
        7'd78: vec_data_084 = data_d1[623:616];
        7'd79: vec_data_084 = data_d1[631:624];
        7'd80: vec_data_084 = data_d1[639:632];
        7'd81: vec_data_084 = data_d1[647:640];
        7'd82: vec_data_084 = data_d1[655:648];
        7'd83: vec_data_084 = data_d1[663:656];
        7'd84: vec_data_084 = data_d1[671:664];
        7'd85: vec_data_084 = data_d1[679:672];
    endcase
end

always @(
  vec_sum_085_d1
  or data_d1
  ) begin
    vec_data_085 = 8'b0;
    case(vec_sum_085_d1)
        7'd1: vec_data_085 = data_d1[7:0];
        7'd2: vec_data_085 = data_d1[15:8];
        7'd3: vec_data_085 = data_d1[23:16];
        7'd4: vec_data_085 = data_d1[31:24];
        7'd5: vec_data_085 = data_d1[39:32];
        7'd6: vec_data_085 = data_d1[47:40];
        7'd7: vec_data_085 = data_d1[55:48];
        7'd8: vec_data_085 = data_d1[63:56];
        7'd9: vec_data_085 = data_d1[71:64];
        7'd10: vec_data_085 = data_d1[79:72];
        7'd11: vec_data_085 = data_d1[87:80];
        7'd12: vec_data_085 = data_d1[95:88];
        7'd13: vec_data_085 = data_d1[103:96];
        7'd14: vec_data_085 = data_d1[111:104];
        7'd15: vec_data_085 = data_d1[119:112];
        7'd16: vec_data_085 = data_d1[127:120];
        7'd17: vec_data_085 = data_d1[135:128];
        7'd18: vec_data_085 = data_d1[143:136];
        7'd19: vec_data_085 = data_d1[151:144];
        7'd20: vec_data_085 = data_d1[159:152];
        7'd21: vec_data_085 = data_d1[167:160];
        7'd22: vec_data_085 = data_d1[175:168];
        7'd23: vec_data_085 = data_d1[183:176];
        7'd24: vec_data_085 = data_d1[191:184];
        7'd25: vec_data_085 = data_d1[199:192];
        7'd26: vec_data_085 = data_d1[207:200];
        7'd27: vec_data_085 = data_d1[215:208];
        7'd28: vec_data_085 = data_d1[223:216];
        7'd29: vec_data_085 = data_d1[231:224];
        7'd30: vec_data_085 = data_d1[239:232];
        7'd31: vec_data_085 = data_d1[247:240];
        7'd32: vec_data_085 = data_d1[255:248];
        7'd33: vec_data_085 = data_d1[263:256];
        7'd34: vec_data_085 = data_d1[271:264];
        7'd35: vec_data_085 = data_d1[279:272];
        7'd36: vec_data_085 = data_d1[287:280];
        7'd37: vec_data_085 = data_d1[295:288];
        7'd38: vec_data_085 = data_d1[303:296];
        7'd39: vec_data_085 = data_d1[311:304];
        7'd40: vec_data_085 = data_d1[319:312];
        7'd41: vec_data_085 = data_d1[327:320];
        7'd42: vec_data_085 = data_d1[335:328];
        7'd43: vec_data_085 = data_d1[343:336];
        7'd44: vec_data_085 = data_d1[351:344];
        7'd45: vec_data_085 = data_d1[359:352];
        7'd46: vec_data_085 = data_d1[367:360];
        7'd47: vec_data_085 = data_d1[375:368];
        7'd48: vec_data_085 = data_d1[383:376];
        7'd49: vec_data_085 = data_d1[391:384];
        7'd50: vec_data_085 = data_d1[399:392];
        7'd51: vec_data_085 = data_d1[407:400];
        7'd52: vec_data_085 = data_d1[415:408];
        7'd53: vec_data_085 = data_d1[423:416];
        7'd54: vec_data_085 = data_d1[431:424];
        7'd55: vec_data_085 = data_d1[439:432];
        7'd56: vec_data_085 = data_d1[447:440];
        7'd57: vec_data_085 = data_d1[455:448];
        7'd58: vec_data_085 = data_d1[463:456];
        7'd59: vec_data_085 = data_d1[471:464];
        7'd60: vec_data_085 = data_d1[479:472];
        7'd61: vec_data_085 = data_d1[487:480];
        7'd62: vec_data_085 = data_d1[495:488];
        7'd63: vec_data_085 = data_d1[503:496];
        7'd64: vec_data_085 = data_d1[511:504];
        7'd65: vec_data_085 = data_d1[519:512];
        7'd66: vec_data_085 = data_d1[527:520];
        7'd67: vec_data_085 = data_d1[535:528];
        7'd68: vec_data_085 = data_d1[543:536];
        7'd69: vec_data_085 = data_d1[551:544];
        7'd70: vec_data_085 = data_d1[559:552];
        7'd71: vec_data_085 = data_d1[567:560];
        7'd72: vec_data_085 = data_d1[575:568];
        7'd73: vec_data_085 = data_d1[583:576];
        7'd74: vec_data_085 = data_d1[591:584];
        7'd75: vec_data_085 = data_d1[599:592];
        7'd76: vec_data_085 = data_d1[607:600];
        7'd77: vec_data_085 = data_d1[615:608];
        7'd78: vec_data_085 = data_d1[623:616];
        7'd79: vec_data_085 = data_d1[631:624];
        7'd80: vec_data_085 = data_d1[639:632];
        7'd81: vec_data_085 = data_d1[647:640];
        7'd82: vec_data_085 = data_d1[655:648];
        7'd83: vec_data_085 = data_d1[663:656];
        7'd84: vec_data_085 = data_d1[671:664];
        7'd85: vec_data_085 = data_d1[679:672];
        7'd86: vec_data_085 = data_d1[687:680];
    endcase
end

always @(
  vec_sum_086_d1
  or data_d1
  ) begin
    vec_data_086 = 8'b0;
    case(vec_sum_086_d1)
        7'd1: vec_data_086 = data_d1[7:0];
        7'd2: vec_data_086 = data_d1[15:8];
        7'd3: vec_data_086 = data_d1[23:16];
        7'd4: vec_data_086 = data_d1[31:24];
        7'd5: vec_data_086 = data_d1[39:32];
        7'd6: vec_data_086 = data_d1[47:40];
        7'd7: vec_data_086 = data_d1[55:48];
        7'd8: vec_data_086 = data_d1[63:56];
        7'd9: vec_data_086 = data_d1[71:64];
        7'd10: vec_data_086 = data_d1[79:72];
        7'd11: vec_data_086 = data_d1[87:80];
        7'd12: vec_data_086 = data_d1[95:88];
        7'd13: vec_data_086 = data_d1[103:96];
        7'd14: vec_data_086 = data_d1[111:104];
        7'd15: vec_data_086 = data_d1[119:112];
        7'd16: vec_data_086 = data_d1[127:120];
        7'd17: vec_data_086 = data_d1[135:128];
        7'd18: vec_data_086 = data_d1[143:136];
        7'd19: vec_data_086 = data_d1[151:144];
        7'd20: vec_data_086 = data_d1[159:152];
        7'd21: vec_data_086 = data_d1[167:160];
        7'd22: vec_data_086 = data_d1[175:168];
        7'd23: vec_data_086 = data_d1[183:176];
        7'd24: vec_data_086 = data_d1[191:184];
        7'd25: vec_data_086 = data_d1[199:192];
        7'd26: vec_data_086 = data_d1[207:200];
        7'd27: vec_data_086 = data_d1[215:208];
        7'd28: vec_data_086 = data_d1[223:216];
        7'd29: vec_data_086 = data_d1[231:224];
        7'd30: vec_data_086 = data_d1[239:232];
        7'd31: vec_data_086 = data_d1[247:240];
        7'd32: vec_data_086 = data_d1[255:248];
        7'd33: vec_data_086 = data_d1[263:256];
        7'd34: vec_data_086 = data_d1[271:264];
        7'd35: vec_data_086 = data_d1[279:272];
        7'd36: vec_data_086 = data_d1[287:280];
        7'd37: vec_data_086 = data_d1[295:288];
        7'd38: vec_data_086 = data_d1[303:296];
        7'd39: vec_data_086 = data_d1[311:304];
        7'd40: vec_data_086 = data_d1[319:312];
        7'd41: vec_data_086 = data_d1[327:320];
        7'd42: vec_data_086 = data_d1[335:328];
        7'd43: vec_data_086 = data_d1[343:336];
        7'd44: vec_data_086 = data_d1[351:344];
        7'd45: vec_data_086 = data_d1[359:352];
        7'd46: vec_data_086 = data_d1[367:360];
        7'd47: vec_data_086 = data_d1[375:368];
        7'd48: vec_data_086 = data_d1[383:376];
        7'd49: vec_data_086 = data_d1[391:384];
        7'd50: vec_data_086 = data_d1[399:392];
        7'd51: vec_data_086 = data_d1[407:400];
        7'd52: vec_data_086 = data_d1[415:408];
        7'd53: vec_data_086 = data_d1[423:416];
        7'd54: vec_data_086 = data_d1[431:424];
        7'd55: vec_data_086 = data_d1[439:432];
        7'd56: vec_data_086 = data_d1[447:440];
        7'd57: vec_data_086 = data_d1[455:448];
        7'd58: vec_data_086 = data_d1[463:456];
        7'd59: vec_data_086 = data_d1[471:464];
        7'd60: vec_data_086 = data_d1[479:472];
        7'd61: vec_data_086 = data_d1[487:480];
        7'd62: vec_data_086 = data_d1[495:488];
        7'd63: vec_data_086 = data_d1[503:496];
        7'd64: vec_data_086 = data_d1[511:504];
        7'd65: vec_data_086 = data_d1[519:512];
        7'd66: vec_data_086 = data_d1[527:520];
        7'd67: vec_data_086 = data_d1[535:528];
        7'd68: vec_data_086 = data_d1[543:536];
        7'd69: vec_data_086 = data_d1[551:544];
        7'd70: vec_data_086 = data_d1[559:552];
        7'd71: vec_data_086 = data_d1[567:560];
        7'd72: vec_data_086 = data_d1[575:568];
        7'd73: vec_data_086 = data_d1[583:576];
        7'd74: vec_data_086 = data_d1[591:584];
        7'd75: vec_data_086 = data_d1[599:592];
        7'd76: vec_data_086 = data_d1[607:600];
        7'd77: vec_data_086 = data_d1[615:608];
        7'd78: vec_data_086 = data_d1[623:616];
        7'd79: vec_data_086 = data_d1[631:624];
        7'd80: vec_data_086 = data_d1[639:632];
        7'd81: vec_data_086 = data_d1[647:640];
        7'd82: vec_data_086 = data_d1[655:648];
        7'd83: vec_data_086 = data_d1[663:656];
        7'd84: vec_data_086 = data_d1[671:664];
        7'd85: vec_data_086 = data_d1[679:672];
        7'd86: vec_data_086 = data_d1[687:680];
        7'd87: vec_data_086 = data_d1[695:688];
    endcase
end

always @(
  vec_sum_087_d1
  or data_d1
  ) begin
    vec_data_087 = 8'b0;
    case(vec_sum_087_d1)
        7'd1: vec_data_087 = data_d1[7:0];
        7'd2: vec_data_087 = data_d1[15:8];
        7'd3: vec_data_087 = data_d1[23:16];
        7'd4: vec_data_087 = data_d1[31:24];
        7'd5: vec_data_087 = data_d1[39:32];
        7'd6: vec_data_087 = data_d1[47:40];
        7'd7: vec_data_087 = data_d1[55:48];
        7'd8: vec_data_087 = data_d1[63:56];
        7'd9: vec_data_087 = data_d1[71:64];
        7'd10: vec_data_087 = data_d1[79:72];
        7'd11: vec_data_087 = data_d1[87:80];
        7'd12: vec_data_087 = data_d1[95:88];
        7'd13: vec_data_087 = data_d1[103:96];
        7'd14: vec_data_087 = data_d1[111:104];
        7'd15: vec_data_087 = data_d1[119:112];
        7'd16: vec_data_087 = data_d1[127:120];
        7'd17: vec_data_087 = data_d1[135:128];
        7'd18: vec_data_087 = data_d1[143:136];
        7'd19: vec_data_087 = data_d1[151:144];
        7'd20: vec_data_087 = data_d1[159:152];
        7'd21: vec_data_087 = data_d1[167:160];
        7'd22: vec_data_087 = data_d1[175:168];
        7'd23: vec_data_087 = data_d1[183:176];
        7'd24: vec_data_087 = data_d1[191:184];
        7'd25: vec_data_087 = data_d1[199:192];
        7'd26: vec_data_087 = data_d1[207:200];
        7'd27: vec_data_087 = data_d1[215:208];
        7'd28: vec_data_087 = data_d1[223:216];
        7'd29: vec_data_087 = data_d1[231:224];
        7'd30: vec_data_087 = data_d1[239:232];
        7'd31: vec_data_087 = data_d1[247:240];
        7'd32: vec_data_087 = data_d1[255:248];
        7'd33: vec_data_087 = data_d1[263:256];
        7'd34: vec_data_087 = data_d1[271:264];
        7'd35: vec_data_087 = data_d1[279:272];
        7'd36: vec_data_087 = data_d1[287:280];
        7'd37: vec_data_087 = data_d1[295:288];
        7'd38: vec_data_087 = data_d1[303:296];
        7'd39: vec_data_087 = data_d1[311:304];
        7'd40: vec_data_087 = data_d1[319:312];
        7'd41: vec_data_087 = data_d1[327:320];
        7'd42: vec_data_087 = data_d1[335:328];
        7'd43: vec_data_087 = data_d1[343:336];
        7'd44: vec_data_087 = data_d1[351:344];
        7'd45: vec_data_087 = data_d1[359:352];
        7'd46: vec_data_087 = data_d1[367:360];
        7'd47: vec_data_087 = data_d1[375:368];
        7'd48: vec_data_087 = data_d1[383:376];
        7'd49: vec_data_087 = data_d1[391:384];
        7'd50: vec_data_087 = data_d1[399:392];
        7'd51: vec_data_087 = data_d1[407:400];
        7'd52: vec_data_087 = data_d1[415:408];
        7'd53: vec_data_087 = data_d1[423:416];
        7'd54: vec_data_087 = data_d1[431:424];
        7'd55: vec_data_087 = data_d1[439:432];
        7'd56: vec_data_087 = data_d1[447:440];
        7'd57: vec_data_087 = data_d1[455:448];
        7'd58: vec_data_087 = data_d1[463:456];
        7'd59: vec_data_087 = data_d1[471:464];
        7'd60: vec_data_087 = data_d1[479:472];
        7'd61: vec_data_087 = data_d1[487:480];
        7'd62: vec_data_087 = data_d1[495:488];
        7'd63: vec_data_087 = data_d1[503:496];
        7'd64: vec_data_087 = data_d1[511:504];
        7'd65: vec_data_087 = data_d1[519:512];
        7'd66: vec_data_087 = data_d1[527:520];
        7'd67: vec_data_087 = data_d1[535:528];
        7'd68: vec_data_087 = data_d1[543:536];
        7'd69: vec_data_087 = data_d1[551:544];
        7'd70: vec_data_087 = data_d1[559:552];
        7'd71: vec_data_087 = data_d1[567:560];
        7'd72: vec_data_087 = data_d1[575:568];
        7'd73: vec_data_087 = data_d1[583:576];
        7'd74: vec_data_087 = data_d1[591:584];
        7'd75: vec_data_087 = data_d1[599:592];
        7'd76: vec_data_087 = data_d1[607:600];
        7'd77: vec_data_087 = data_d1[615:608];
        7'd78: vec_data_087 = data_d1[623:616];
        7'd79: vec_data_087 = data_d1[631:624];
        7'd80: vec_data_087 = data_d1[639:632];
        7'd81: vec_data_087 = data_d1[647:640];
        7'd82: vec_data_087 = data_d1[655:648];
        7'd83: vec_data_087 = data_d1[663:656];
        7'd84: vec_data_087 = data_d1[671:664];
        7'd85: vec_data_087 = data_d1[679:672];
        7'd86: vec_data_087 = data_d1[687:680];
        7'd87: vec_data_087 = data_d1[695:688];
        7'd88: vec_data_087 = data_d1[703:696];
    endcase
end

always @(
  vec_sum_088_d1
  or data_d1
  ) begin
    vec_data_088 = 8'b0;
    case(vec_sum_088_d1)
        7'd1: vec_data_088 = data_d1[7:0];
        7'd2: vec_data_088 = data_d1[15:8];
        7'd3: vec_data_088 = data_d1[23:16];
        7'd4: vec_data_088 = data_d1[31:24];
        7'd5: vec_data_088 = data_d1[39:32];
        7'd6: vec_data_088 = data_d1[47:40];
        7'd7: vec_data_088 = data_d1[55:48];
        7'd8: vec_data_088 = data_d1[63:56];
        7'd9: vec_data_088 = data_d1[71:64];
        7'd10: vec_data_088 = data_d1[79:72];
        7'd11: vec_data_088 = data_d1[87:80];
        7'd12: vec_data_088 = data_d1[95:88];
        7'd13: vec_data_088 = data_d1[103:96];
        7'd14: vec_data_088 = data_d1[111:104];
        7'd15: vec_data_088 = data_d1[119:112];
        7'd16: vec_data_088 = data_d1[127:120];
        7'd17: vec_data_088 = data_d1[135:128];
        7'd18: vec_data_088 = data_d1[143:136];
        7'd19: vec_data_088 = data_d1[151:144];
        7'd20: vec_data_088 = data_d1[159:152];
        7'd21: vec_data_088 = data_d1[167:160];
        7'd22: vec_data_088 = data_d1[175:168];
        7'd23: vec_data_088 = data_d1[183:176];
        7'd24: vec_data_088 = data_d1[191:184];
        7'd25: vec_data_088 = data_d1[199:192];
        7'd26: vec_data_088 = data_d1[207:200];
        7'd27: vec_data_088 = data_d1[215:208];
        7'd28: vec_data_088 = data_d1[223:216];
        7'd29: vec_data_088 = data_d1[231:224];
        7'd30: vec_data_088 = data_d1[239:232];
        7'd31: vec_data_088 = data_d1[247:240];
        7'd32: vec_data_088 = data_d1[255:248];
        7'd33: vec_data_088 = data_d1[263:256];
        7'd34: vec_data_088 = data_d1[271:264];
        7'd35: vec_data_088 = data_d1[279:272];
        7'd36: vec_data_088 = data_d1[287:280];
        7'd37: vec_data_088 = data_d1[295:288];
        7'd38: vec_data_088 = data_d1[303:296];
        7'd39: vec_data_088 = data_d1[311:304];
        7'd40: vec_data_088 = data_d1[319:312];
        7'd41: vec_data_088 = data_d1[327:320];
        7'd42: vec_data_088 = data_d1[335:328];
        7'd43: vec_data_088 = data_d1[343:336];
        7'd44: vec_data_088 = data_d1[351:344];
        7'd45: vec_data_088 = data_d1[359:352];
        7'd46: vec_data_088 = data_d1[367:360];
        7'd47: vec_data_088 = data_d1[375:368];
        7'd48: vec_data_088 = data_d1[383:376];
        7'd49: vec_data_088 = data_d1[391:384];
        7'd50: vec_data_088 = data_d1[399:392];
        7'd51: vec_data_088 = data_d1[407:400];
        7'd52: vec_data_088 = data_d1[415:408];
        7'd53: vec_data_088 = data_d1[423:416];
        7'd54: vec_data_088 = data_d1[431:424];
        7'd55: vec_data_088 = data_d1[439:432];
        7'd56: vec_data_088 = data_d1[447:440];
        7'd57: vec_data_088 = data_d1[455:448];
        7'd58: vec_data_088 = data_d1[463:456];
        7'd59: vec_data_088 = data_d1[471:464];
        7'd60: vec_data_088 = data_d1[479:472];
        7'd61: vec_data_088 = data_d1[487:480];
        7'd62: vec_data_088 = data_d1[495:488];
        7'd63: vec_data_088 = data_d1[503:496];
        7'd64: vec_data_088 = data_d1[511:504];
        7'd65: vec_data_088 = data_d1[519:512];
        7'd66: vec_data_088 = data_d1[527:520];
        7'd67: vec_data_088 = data_d1[535:528];
        7'd68: vec_data_088 = data_d1[543:536];
        7'd69: vec_data_088 = data_d1[551:544];
        7'd70: vec_data_088 = data_d1[559:552];
        7'd71: vec_data_088 = data_d1[567:560];
        7'd72: vec_data_088 = data_d1[575:568];
        7'd73: vec_data_088 = data_d1[583:576];
        7'd74: vec_data_088 = data_d1[591:584];
        7'd75: vec_data_088 = data_d1[599:592];
        7'd76: vec_data_088 = data_d1[607:600];
        7'd77: vec_data_088 = data_d1[615:608];
        7'd78: vec_data_088 = data_d1[623:616];
        7'd79: vec_data_088 = data_d1[631:624];
        7'd80: vec_data_088 = data_d1[639:632];
        7'd81: vec_data_088 = data_d1[647:640];
        7'd82: vec_data_088 = data_d1[655:648];
        7'd83: vec_data_088 = data_d1[663:656];
        7'd84: vec_data_088 = data_d1[671:664];
        7'd85: vec_data_088 = data_d1[679:672];
        7'd86: vec_data_088 = data_d1[687:680];
        7'd87: vec_data_088 = data_d1[695:688];
        7'd88: vec_data_088 = data_d1[703:696];
        7'd89: vec_data_088 = data_d1[711:704];
    endcase
end

always @(
  vec_sum_089_d1
  or data_d1
  ) begin
    vec_data_089 = 8'b0;
    case(vec_sum_089_d1)
        7'd1: vec_data_089 = data_d1[7:0];
        7'd2: vec_data_089 = data_d1[15:8];
        7'd3: vec_data_089 = data_d1[23:16];
        7'd4: vec_data_089 = data_d1[31:24];
        7'd5: vec_data_089 = data_d1[39:32];
        7'd6: vec_data_089 = data_d1[47:40];
        7'd7: vec_data_089 = data_d1[55:48];
        7'd8: vec_data_089 = data_d1[63:56];
        7'd9: vec_data_089 = data_d1[71:64];
        7'd10: vec_data_089 = data_d1[79:72];
        7'd11: vec_data_089 = data_d1[87:80];
        7'd12: vec_data_089 = data_d1[95:88];
        7'd13: vec_data_089 = data_d1[103:96];
        7'd14: vec_data_089 = data_d1[111:104];
        7'd15: vec_data_089 = data_d1[119:112];
        7'd16: vec_data_089 = data_d1[127:120];
        7'd17: vec_data_089 = data_d1[135:128];
        7'd18: vec_data_089 = data_d1[143:136];
        7'd19: vec_data_089 = data_d1[151:144];
        7'd20: vec_data_089 = data_d1[159:152];
        7'd21: vec_data_089 = data_d1[167:160];
        7'd22: vec_data_089 = data_d1[175:168];
        7'd23: vec_data_089 = data_d1[183:176];
        7'd24: vec_data_089 = data_d1[191:184];
        7'd25: vec_data_089 = data_d1[199:192];
        7'd26: vec_data_089 = data_d1[207:200];
        7'd27: vec_data_089 = data_d1[215:208];
        7'd28: vec_data_089 = data_d1[223:216];
        7'd29: vec_data_089 = data_d1[231:224];
        7'd30: vec_data_089 = data_d1[239:232];
        7'd31: vec_data_089 = data_d1[247:240];
        7'd32: vec_data_089 = data_d1[255:248];
        7'd33: vec_data_089 = data_d1[263:256];
        7'd34: vec_data_089 = data_d1[271:264];
        7'd35: vec_data_089 = data_d1[279:272];
        7'd36: vec_data_089 = data_d1[287:280];
        7'd37: vec_data_089 = data_d1[295:288];
        7'd38: vec_data_089 = data_d1[303:296];
        7'd39: vec_data_089 = data_d1[311:304];
        7'd40: vec_data_089 = data_d1[319:312];
        7'd41: vec_data_089 = data_d1[327:320];
        7'd42: vec_data_089 = data_d1[335:328];
        7'd43: vec_data_089 = data_d1[343:336];
        7'd44: vec_data_089 = data_d1[351:344];
        7'd45: vec_data_089 = data_d1[359:352];
        7'd46: vec_data_089 = data_d1[367:360];
        7'd47: vec_data_089 = data_d1[375:368];
        7'd48: vec_data_089 = data_d1[383:376];
        7'd49: vec_data_089 = data_d1[391:384];
        7'd50: vec_data_089 = data_d1[399:392];
        7'd51: vec_data_089 = data_d1[407:400];
        7'd52: vec_data_089 = data_d1[415:408];
        7'd53: vec_data_089 = data_d1[423:416];
        7'd54: vec_data_089 = data_d1[431:424];
        7'd55: vec_data_089 = data_d1[439:432];
        7'd56: vec_data_089 = data_d1[447:440];
        7'd57: vec_data_089 = data_d1[455:448];
        7'd58: vec_data_089 = data_d1[463:456];
        7'd59: vec_data_089 = data_d1[471:464];
        7'd60: vec_data_089 = data_d1[479:472];
        7'd61: vec_data_089 = data_d1[487:480];
        7'd62: vec_data_089 = data_d1[495:488];
        7'd63: vec_data_089 = data_d1[503:496];
        7'd64: vec_data_089 = data_d1[511:504];
        7'd65: vec_data_089 = data_d1[519:512];
        7'd66: vec_data_089 = data_d1[527:520];
        7'd67: vec_data_089 = data_d1[535:528];
        7'd68: vec_data_089 = data_d1[543:536];
        7'd69: vec_data_089 = data_d1[551:544];
        7'd70: vec_data_089 = data_d1[559:552];
        7'd71: vec_data_089 = data_d1[567:560];
        7'd72: vec_data_089 = data_d1[575:568];
        7'd73: vec_data_089 = data_d1[583:576];
        7'd74: vec_data_089 = data_d1[591:584];
        7'd75: vec_data_089 = data_d1[599:592];
        7'd76: vec_data_089 = data_d1[607:600];
        7'd77: vec_data_089 = data_d1[615:608];
        7'd78: vec_data_089 = data_d1[623:616];
        7'd79: vec_data_089 = data_d1[631:624];
        7'd80: vec_data_089 = data_d1[639:632];
        7'd81: vec_data_089 = data_d1[647:640];
        7'd82: vec_data_089 = data_d1[655:648];
        7'd83: vec_data_089 = data_d1[663:656];
        7'd84: vec_data_089 = data_d1[671:664];
        7'd85: vec_data_089 = data_d1[679:672];
        7'd86: vec_data_089 = data_d1[687:680];
        7'd87: vec_data_089 = data_d1[695:688];
        7'd88: vec_data_089 = data_d1[703:696];
        7'd89: vec_data_089 = data_d1[711:704];
        7'd90: vec_data_089 = data_d1[719:712];
    endcase
end

always @(
  vec_sum_090_d1
  or data_d1
  ) begin
    vec_data_090 = 8'b0;
    case(vec_sum_090_d1)
        7'd1: vec_data_090 = data_d1[7:0];
        7'd2: vec_data_090 = data_d1[15:8];
        7'd3: vec_data_090 = data_d1[23:16];
        7'd4: vec_data_090 = data_d1[31:24];
        7'd5: vec_data_090 = data_d1[39:32];
        7'd6: vec_data_090 = data_d1[47:40];
        7'd7: vec_data_090 = data_d1[55:48];
        7'd8: vec_data_090 = data_d1[63:56];
        7'd9: vec_data_090 = data_d1[71:64];
        7'd10: vec_data_090 = data_d1[79:72];
        7'd11: vec_data_090 = data_d1[87:80];
        7'd12: vec_data_090 = data_d1[95:88];
        7'd13: vec_data_090 = data_d1[103:96];
        7'd14: vec_data_090 = data_d1[111:104];
        7'd15: vec_data_090 = data_d1[119:112];
        7'd16: vec_data_090 = data_d1[127:120];
        7'd17: vec_data_090 = data_d1[135:128];
        7'd18: vec_data_090 = data_d1[143:136];
        7'd19: vec_data_090 = data_d1[151:144];
        7'd20: vec_data_090 = data_d1[159:152];
        7'd21: vec_data_090 = data_d1[167:160];
        7'd22: vec_data_090 = data_d1[175:168];
        7'd23: vec_data_090 = data_d1[183:176];
        7'd24: vec_data_090 = data_d1[191:184];
        7'd25: vec_data_090 = data_d1[199:192];
        7'd26: vec_data_090 = data_d1[207:200];
        7'd27: vec_data_090 = data_d1[215:208];
        7'd28: vec_data_090 = data_d1[223:216];
        7'd29: vec_data_090 = data_d1[231:224];
        7'd30: vec_data_090 = data_d1[239:232];
        7'd31: vec_data_090 = data_d1[247:240];
        7'd32: vec_data_090 = data_d1[255:248];
        7'd33: vec_data_090 = data_d1[263:256];
        7'd34: vec_data_090 = data_d1[271:264];
        7'd35: vec_data_090 = data_d1[279:272];
        7'd36: vec_data_090 = data_d1[287:280];
        7'd37: vec_data_090 = data_d1[295:288];
        7'd38: vec_data_090 = data_d1[303:296];
        7'd39: vec_data_090 = data_d1[311:304];
        7'd40: vec_data_090 = data_d1[319:312];
        7'd41: vec_data_090 = data_d1[327:320];
        7'd42: vec_data_090 = data_d1[335:328];
        7'd43: vec_data_090 = data_d1[343:336];
        7'd44: vec_data_090 = data_d1[351:344];
        7'd45: vec_data_090 = data_d1[359:352];
        7'd46: vec_data_090 = data_d1[367:360];
        7'd47: vec_data_090 = data_d1[375:368];
        7'd48: vec_data_090 = data_d1[383:376];
        7'd49: vec_data_090 = data_d1[391:384];
        7'd50: vec_data_090 = data_d1[399:392];
        7'd51: vec_data_090 = data_d1[407:400];
        7'd52: vec_data_090 = data_d1[415:408];
        7'd53: vec_data_090 = data_d1[423:416];
        7'd54: vec_data_090 = data_d1[431:424];
        7'd55: vec_data_090 = data_d1[439:432];
        7'd56: vec_data_090 = data_d1[447:440];
        7'd57: vec_data_090 = data_d1[455:448];
        7'd58: vec_data_090 = data_d1[463:456];
        7'd59: vec_data_090 = data_d1[471:464];
        7'd60: vec_data_090 = data_d1[479:472];
        7'd61: vec_data_090 = data_d1[487:480];
        7'd62: vec_data_090 = data_d1[495:488];
        7'd63: vec_data_090 = data_d1[503:496];
        7'd64: vec_data_090 = data_d1[511:504];
        7'd65: vec_data_090 = data_d1[519:512];
        7'd66: vec_data_090 = data_d1[527:520];
        7'd67: vec_data_090 = data_d1[535:528];
        7'd68: vec_data_090 = data_d1[543:536];
        7'd69: vec_data_090 = data_d1[551:544];
        7'd70: vec_data_090 = data_d1[559:552];
        7'd71: vec_data_090 = data_d1[567:560];
        7'd72: vec_data_090 = data_d1[575:568];
        7'd73: vec_data_090 = data_d1[583:576];
        7'd74: vec_data_090 = data_d1[591:584];
        7'd75: vec_data_090 = data_d1[599:592];
        7'd76: vec_data_090 = data_d1[607:600];
        7'd77: vec_data_090 = data_d1[615:608];
        7'd78: vec_data_090 = data_d1[623:616];
        7'd79: vec_data_090 = data_d1[631:624];
        7'd80: vec_data_090 = data_d1[639:632];
        7'd81: vec_data_090 = data_d1[647:640];
        7'd82: vec_data_090 = data_d1[655:648];
        7'd83: vec_data_090 = data_d1[663:656];
        7'd84: vec_data_090 = data_d1[671:664];
        7'd85: vec_data_090 = data_d1[679:672];
        7'd86: vec_data_090 = data_d1[687:680];
        7'd87: vec_data_090 = data_d1[695:688];
        7'd88: vec_data_090 = data_d1[703:696];
        7'd89: vec_data_090 = data_d1[711:704];
        7'd90: vec_data_090 = data_d1[719:712];
        7'd91: vec_data_090 = data_d1[727:720];
    endcase
end

always @(
  vec_sum_091_d1
  or data_d1
  ) begin
    vec_data_091 = 8'b0;
    case(vec_sum_091_d1)
        7'd1: vec_data_091 = data_d1[7:0];
        7'd2: vec_data_091 = data_d1[15:8];
        7'd3: vec_data_091 = data_d1[23:16];
        7'd4: vec_data_091 = data_d1[31:24];
        7'd5: vec_data_091 = data_d1[39:32];
        7'd6: vec_data_091 = data_d1[47:40];
        7'd7: vec_data_091 = data_d1[55:48];
        7'd8: vec_data_091 = data_d1[63:56];
        7'd9: vec_data_091 = data_d1[71:64];
        7'd10: vec_data_091 = data_d1[79:72];
        7'd11: vec_data_091 = data_d1[87:80];
        7'd12: vec_data_091 = data_d1[95:88];
        7'd13: vec_data_091 = data_d1[103:96];
        7'd14: vec_data_091 = data_d1[111:104];
        7'd15: vec_data_091 = data_d1[119:112];
        7'd16: vec_data_091 = data_d1[127:120];
        7'd17: vec_data_091 = data_d1[135:128];
        7'd18: vec_data_091 = data_d1[143:136];
        7'd19: vec_data_091 = data_d1[151:144];
        7'd20: vec_data_091 = data_d1[159:152];
        7'd21: vec_data_091 = data_d1[167:160];
        7'd22: vec_data_091 = data_d1[175:168];
        7'd23: vec_data_091 = data_d1[183:176];
        7'd24: vec_data_091 = data_d1[191:184];
        7'd25: vec_data_091 = data_d1[199:192];
        7'd26: vec_data_091 = data_d1[207:200];
        7'd27: vec_data_091 = data_d1[215:208];
        7'd28: vec_data_091 = data_d1[223:216];
        7'd29: vec_data_091 = data_d1[231:224];
        7'd30: vec_data_091 = data_d1[239:232];
        7'd31: vec_data_091 = data_d1[247:240];
        7'd32: vec_data_091 = data_d1[255:248];
        7'd33: vec_data_091 = data_d1[263:256];
        7'd34: vec_data_091 = data_d1[271:264];
        7'd35: vec_data_091 = data_d1[279:272];
        7'd36: vec_data_091 = data_d1[287:280];
        7'd37: vec_data_091 = data_d1[295:288];
        7'd38: vec_data_091 = data_d1[303:296];
        7'd39: vec_data_091 = data_d1[311:304];
        7'd40: vec_data_091 = data_d1[319:312];
        7'd41: vec_data_091 = data_d1[327:320];
        7'd42: vec_data_091 = data_d1[335:328];
        7'd43: vec_data_091 = data_d1[343:336];
        7'd44: vec_data_091 = data_d1[351:344];
        7'd45: vec_data_091 = data_d1[359:352];
        7'd46: vec_data_091 = data_d1[367:360];
        7'd47: vec_data_091 = data_d1[375:368];
        7'd48: vec_data_091 = data_d1[383:376];
        7'd49: vec_data_091 = data_d1[391:384];
        7'd50: vec_data_091 = data_d1[399:392];
        7'd51: vec_data_091 = data_d1[407:400];
        7'd52: vec_data_091 = data_d1[415:408];
        7'd53: vec_data_091 = data_d1[423:416];
        7'd54: vec_data_091 = data_d1[431:424];
        7'd55: vec_data_091 = data_d1[439:432];
        7'd56: vec_data_091 = data_d1[447:440];
        7'd57: vec_data_091 = data_d1[455:448];
        7'd58: vec_data_091 = data_d1[463:456];
        7'd59: vec_data_091 = data_d1[471:464];
        7'd60: vec_data_091 = data_d1[479:472];
        7'd61: vec_data_091 = data_d1[487:480];
        7'd62: vec_data_091 = data_d1[495:488];
        7'd63: vec_data_091 = data_d1[503:496];
        7'd64: vec_data_091 = data_d1[511:504];
        7'd65: vec_data_091 = data_d1[519:512];
        7'd66: vec_data_091 = data_d1[527:520];
        7'd67: vec_data_091 = data_d1[535:528];
        7'd68: vec_data_091 = data_d1[543:536];
        7'd69: vec_data_091 = data_d1[551:544];
        7'd70: vec_data_091 = data_d1[559:552];
        7'd71: vec_data_091 = data_d1[567:560];
        7'd72: vec_data_091 = data_d1[575:568];
        7'd73: vec_data_091 = data_d1[583:576];
        7'd74: vec_data_091 = data_d1[591:584];
        7'd75: vec_data_091 = data_d1[599:592];
        7'd76: vec_data_091 = data_d1[607:600];
        7'd77: vec_data_091 = data_d1[615:608];
        7'd78: vec_data_091 = data_d1[623:616];
        7'd79: vec_data_091 = data_d1[631:624];
        7'd80: vec_data_091 = data_d1[639:632];
        7'd81: vec_data_091 = data_d1[647:640];
        7'd82: vec_data_091 = data_d1[655:648];
        7'd83: vec_data_091 = data_d1[663:656];
        7'd84: vec_data_091 = data_d1[671:664];
        7'd85: vec_data_091 = data_d1[679:672];
        7'd86: vec_data_091 = data_d1[687:680];
        7'd87: vec_data_091 = data_d1[695:688];
        7'd88: vec_data_091 = data_d1[703:696];
        7'd89: vec_data_091 = data_d1[711:704];
        7'd90: vec_data_091 = data_d1[719:712];
        7'd91: vec_data_091 = data_d1[727:720];
        7'd92: vec_data_091 = data_d1[735:728];
    endcase
end

always @(
  vec_sum_092_d1
  or data_d1
  ) begin
    vec_data_092 = 8'b0;
    case(vec_sum_092_d1)
        7'd1: vec_data_092 = data_d1[7:0];
        7'd2: vec_data_092 = data_d1[15:8];
        7'd3: vec_data_092 = data_d1[23:16];
        7'd4: vec_data_092 = data_d1[31:24];
        7'd5: vec_data_092 = data_d1[39:32];
        7'd6: vec_data_092 = data_d1[47:40];
        7'd7: vec_data_092 = data_d1[55:48];
        7'd8: vec_data_092 = data_d1[63:56];
        7'd9: vec_data_092 = data_d1[71:64];
        7'd10: vec_data_092 = data_d1[79:72];
        7'd11: vec_data_092 = data_d1[87:80];
        7'd12: vec_data_092 = data_d1[95:88];
        7'd13: vec_data_092 = data_d1[103:96];
        7'd14: vec_data_092 = data_d1[111:104];
        7'd15: vec_data_092 = data_d1[119:112];
        7'd16: vec_data_092 = data_d1[127:120];
        7'd17: vec_data_092 = data_d1[135:128];
        7'd18: vec_data_092 = data_d1[143:136];
        7'd19: vec_data_092 = data_d1[151:144];
        7'd20: vec_data_092 = data_d1[159:152];
        7'd21: vec_data_092 = data_d1[167:160];
        7'd22: vec_data_092 = data_d1[175:168];
        7'd23: vec_data_092 = data_d1[183:176];
        7'd24: vec_data_092 = data_d1[191:184];
        7'd25: vec_data_092 = data_d1[199:192];
        7'd26: vec_data_092 = data_d1[207:200];
        7'd27: vec_data_092 = data_d1[215:208];
        7'd28: vec_data_092 = data_d1[223:216];
        7'd29: vec_data_092 = data_d1[231:224];
        7'd30: vec_data_092 = data_d1[239:232];
        7'd31: vec_data_092 = data_d1[247:240];
        7'd32: vec_data_092 = data_d1[255:248];
        7'd33: vec_data_092 = data_d1[263:256];
        7'd34: vec_data_092 = data_d1[271:264];
        7'd35: vec_data_092 = data_d1[279:272];
        7'd36: vec_data_092 = data_d1[287:280];
        7'd37: vec_data_092 = data_d1[295:288];
        7'd38: vec_data_092 = data_d1[303:296];
        7'd39: vec_data_092 = data_d1[311:304];
        7'd40: vec_data_092 = data_d1[319:312];
        7'd41: vec_data_092 = data_d1[327:320];
        7'd42: vec_data_092 = data_d1[335:328];
        7'd43: vec_data_092 = data_d1[343:336];
        7'd44: vec_data_092 = data_d1[351:344];
        7'd45: vec_data_092 = data_d1[359:352];
        7'd46: vec_data_092 = data_d1[367:360];
        7'd47: vec_data_092 = data_d1[375:368];
        7'd48: vec_data_092 = data_d1[383:376];
        7'd49: vec_data_092 = data_d1[391:384];
        7'd50: vec_data_092 = data_d1[399:392];
        7'd51: vec_data_092 = data_d1[407:400];
        7'd52: vec_data_092 = data_d1[415:408];
        7'd53: vec_data_092 = data_d1[423:416];
        7'd54: vec_data_092 = data_d1[431:424];
        7'd55: vec_data_092 = data_d1[439:432];
        7'd56: vec_data_092 = data_d1[447:440];
        7'd57: vec_data_092 = data_d1[455:448];
        7'd58: vec_data_092 = data_d1[463:456];
        7'd59: vec_data_092 = data_d1[471:464];
        7'd60: vec_data_092 = data_d1[479:472];
        7'd61: vec_data_092 = data_d1[487:480];
        7'd62: vec_data_092 = data_d1[495:488];
        7'd63: vec_data_092 = data_d1[503:496];
        7'd64: vec_data_092 = data_d1[511:504];
        7'd65: vec_data_092 = data_d1[519:512];
        7'd66: vec_data_092 = data_d1[527:520];
        7'd67: vec_data_092 = data_d1[535:528];
        7'd68: vec_data_092 = data_d1[543:536];
        7'd69: vec_data_092 = data_d1[551:544];
        7'd70: vec_data_092 = data_d1[559:552];
        7'd71: vec_data_092 = data_d1[567:560];
        7'd72: vec_data_092 = data_d1[575:568];
        7'd73: vec_data_092 = data_d1[583:576];
        7'd74: vec_data_092 = data_d1[591:584];
        7'd75: vec_data_092 = data_d1[599:592];
        7'd76: vec_data_092 = data_d1[607:600];
        7'd77: vec_data_092 = data_d1[615:608];
        7'd78: vec_data_092 = data_d1[623:616];
        7'd79: vec_data_092 = data_d1[631:624];
        7'd80: vec_data_092 = data_d1[639:632];
        7'd81: vec_data_092 = data_d1[647:640];
        7'd82: vec_data_092 = data_d1[655:648];
        7'd83: vec_data_092 = data_d1[663:656];
        7'd84: vec_data_092 = data_d1[671:664];
        7'd85: vec_data_092 = data_d1[679:672];
        7'd86: vec_data_092 = data_d1[687:680];
        7'd87: vec_data_092 = data_d1[695:688];
        7'd88: vec_data_092 = data_d1[703:696];
        7'd89: vec_data_092 = data_d1[711:704];
        7'd90: vec_data_092 = data_d1[719:712];
        7'd91: vec_data_092 = data_d1[727:720];
        7'd92: vec_data_092 = data_d1[735:728];
        7'd93: vec_data_092 = data_d1[743:736];
    endcase
end

always @(
  vec_sum_093_d1
  or data_d1
  ) begin
    vec_data_093 = 8'b0;
    case(vec_sum_093_d1)
        7'd1: vec_data_093 = data_d1[7:0];
        7'd2: vec_data_093 = data_d1[15:8];
        7'd3: vec_data_093 = data_d1[23:16];
        7'd4: vec_data_093 = data_d1[31:24];
        7'd5: vec_data_093 = data_d1[39:32];
        7'd6: vec_data_093 = data_d1[47:40];
        7'd7: vec_data_093 = data_d1[55:48];
        7'd8: vec_data_093 = data_d1[63:56];
        7'd9: vec_data_093 = data_d1[71:64];
        7'd10: vec_data_093 = data_d1[79:72];
        7'd11: vec_data_093 = data_d1[87:80];
        7'd12: vec_data_093 = data_d1[95:88];
        7'd13: vec_data_093 = data_d1[103:96];
        7'd14: vec_data_093 = data_d1[111:104];
        7'd15: vec_data_093 = data_d1[119:112];
        7'd16: vec_data_093 = data_d1[127:120];
        7'd17: vec_data_093 = data_d1[135:128];
        7'd18: vec_data_093 = data_d1[143:136];
        7'd19: vec_data_093 = data_d1[151:144];
        7'd20: vec_data_093 = data_d1[159:152];
        7'd21: vec_data_093 = data_d1[167:160];
        7'd22: vec_data_093 = data_d1[175:168];
        7'd23: vec_data_093 = data_d1[183:176];
        7'd24: vec_data_093 = data_d1[191:184];
        7'd25: vec_data_093 = data_d1[199:192];
        7'd26: vec_data_093 = data_d1[207:200];
        7'd27: vec_data_093 = data_d1[215:208];
        7'd28: vec_data_093 = data_d1[223:216];
        7'd29: vec_data_093 = data_d1[231:224];
        7'd30: vec_data_093 = data_d1[239:232];
        7'd31: vec_data_093 = data_d1[247:240];
        7'd32: vec_data_093 = data_d1[255:248];
        7'd33: vec_data_093 = data_d1[263:256];
        7'd34: vec_data_093 = data_d1[271:264];
        7'd35: vec_data_093 = data_d1[279:272];
        7'd36: vec_data_093 = data_d1[287:280];
        7'd37: vec_data_093 = data_d1[295:288];
        7'd38: vec_data_093 = data_d1[303:296];
        7'd39: vec_data_093 = data_d1[311:304];
        7'd40: vec_data_093 = data_d1[319:312];
        7'd41: vec_data_093 = data_d1[327:320];
        7'd42: vec_data_093 = data_d1[335:328];
        7'd43: vec_data_093 = data_d1[343:336];
        7'd44: vec_data_093 = data_d1[351:344];
        7'd45: vec_data_093 = data_d1[359:352];
        7'd46: vec_data_093 = data_d1[367:360];
        7'd47: vec_data_093 = data_d1[375:368];
        7'd48: vec_data_093 = data_d1[383:376];
        7'd49: vec_data_093 = data_d1[391:384];
        7'd50: vec_data_093 = data_d1[399:392];
        7'd51: vec_data_093 = data_d1[407:400];
        7'd52: vec_data_093 = data_d1[415:408];
        7'd53: vec_data_093 = data_d1[423:416];
        7'd54: vec_data_093 = data_d1[431:424];
        7'd55: vec_data_093 = data_d1[439:432];
        7'd56: vec_data_093 = data_d1[447:440];
        7'd57: vec_data_093 = data_d1[455:448];
        7'd58: vec_data_093 = data_d1[463:456];
        7'd59: vec_data_093 = data_d1[471:464];
        7'd60: vec_data_093 = data_d1[479:472];
        7'd61: vec_data_093 = data_d1[487:480];
        7'd62: vec_data_093 = data_d1[495:488];
        7'd63: vec_data_093 = data_d1[503:496];
        7'd64: vec_data_093 = data_d1[511:504];
        7'd65: vec_data_093 = data_d1[519:512];
        7'd66: vec_data_093 = data_d1[527:520];
        7'd67: vec_data_093 = data_d1[535:528];
        7'd68: vec_data_093 = data_d1[543:536];
        7'd69: vec_data_093 = data_d1[551:544];
        7'd70: vec_data_093 = data_d1[559:552];
        7'd71: vec_data_093 = data_d1[567:560];
        7'd72: vec_data_093 = data_d1[575:568];
        7'd73: vec_data_093 = data_d1[583:576];
        7'd74: vec_data_093 = data_d1[591:584];
        7'd75: vec_data_093 = data_d1[599:592];
        7'd76: vec_data_093 = data_d1[607:600];
        7'd77: vec_data_093 = data_d1[615:608];
        7'd78: vec_data_093 = data_d1[623:616];
        7'd79: vec_data_093 = data_d1[631:624];
        7'd80: vec_data_093 = data_d1[639:632];
        7'd81: vec_data_093 = data_d1[647:640];
        7'd82: vec_data_093 = data_d1[655:648];
        7'd83: vec_data_093 = data_d1[663:656];
        7'd84: vec_data_093 = data_d1[671:664];
        7'd85: vec_data_093 = data_d1[679:672];
        7'd86: vec_data_093 = data_d1[687:680];
        7'd87: vec_data_093 = data_d1[695:688];
        7'd88: vec_data_093 = data_d1[703:696];
        7'd89: vec_data_093 = data_d1[711:704];
        7'd90: vec_data_093 = data_d1[719:712];
        7'd91: vec_data_093 = data_d1[727:720];
        7'd92: vec_data_093 = data_d1[735:728];
        7'd93: vec_data_093 = data_d1[743:736];
        7'd94: vec_data_093 = data_d1[751:744];
    endcase
end

always @(
  vec_sum_094_d1
  or data_d1
  ) begin
    vec_data_094 = 8'b0;
    case(vec_sum_094_d1)
        7'd1: vec_data_094 = data_d1[7:0];
        7'd2: vec_data_094 = data_d1[15:8];
        7'd3: vec_data_094 = data_d1[23:16];
        7'd4: vec_data_094 = data_d1[31:24];
        7'd5: vec_data_094 = data_d1[39:32];
        7'd6: vec_data_094 = data_d1[47:40];
        7'd7: vec_data_094 = data_d1[55:48];
        7'd8: vec_data_094 = data_d1[63:56];
        7'd9: vec_data_094 = data_d1[71:64];
        7'd10: vec_data_094 = data_d1[79:72];
        7'd11: vec_data_094 = data_d1[87:80];
        7'd12: vec_data_094 = data_d1[95:88];
        7'd13: vec_data_094 = data_d1[103:96];
        7'd14: vec_data_094 = data_d1[111:104];
        7'd15: vec_data_094 = data_d1[119:112];
        7'd16: vec_data_094 = data_d1[127:120];
        7'd17: vec_data_094 = data_d1[135:128];
        7'd18: vec_data_094 = data_d1[143:136];
        7'd19: vec_data_094 = data_d1[151:144];
        7'd20: vec_data_094 = data_d1[159:152];
        7'd21: vec_data_094 = data_d1[167:160];
        7'd22: vec_data_094 = data_d1[175:168];
        7'd23: vec_data_094 = data_d1[183:176];
        7'd24: vec_data_094 = data_d1[191:184];
        7'd25: vec_data_094 = data_d1[199:192];
        7'd26: vec_data_094 = data_d1[207:200];
        7'd27: vec_data_094 = data_d1[215:208];
        7'd28: vec_data_094 = data_d1[223:216];
        7'd29: vec_data_094 = data_d1[231:224];
        7'd30: vec_data_094 = data_d1[239:232];
        7'd31: vec_data_094 = data_d1[247:240];
        7'd32: vec_data_094 = data_d1[255:248];
        7'd33: vec_data_094 = data_d1[263:256];
        7'd34: vec_data_094 = data_d1[271:264];
        7'd35: vec_data_094 = data_d1[279:272];
        7'd36: vec_data_094 = data_d1[287:280];
        7'd37: vec_data_094 = data_d1[295:288];
        7'd38: vec_data_094 = data_d1[303:296];
        7'd39: vec_data_094 = data_d1[311:304];
        7'd40: vec_data_094 = data_d1[319:312];
        7'd41: vec_data_094 = data_d1[327:320];
        7'd42: vec_data_094 = data_d1[335:328];
        7'd43: vec_data_094 = data_d1[343:336];
        7'd44: vec_data_094 = data_d1[351:344];
        7'd45: vec_data_094 = data_d1[359:352];
        7'd46: vec_data_094 = data_d1[367:360];
        7'd47: vec_data_094 = data_d1[375:368];
        7'd48: vec_data_094 = data_d1[383:376];
        7'd49: vec_data_094 = data_d1[391:384];
        7'd50: vec_data_094 = data_d1[399:392];
        7'd51: vec_data_094 = data_d1[407:400];
        7'd52: vec_data_094 = data_d1[415:408];
        7'd53: vec_data_094 = data_d1[423:416];
        7'd54: vec_data_094 = data_d1[431:424];
        7'd55: vec_data_094 = data_d1[439:432];
        7'd56: vec_data_094 = data_d1[447:440];
        7'd57: vec_data_094 = data_d1[455:448];
        7'd58: vec_data_094 = data_d1[463:456];
        7'd59: vec_data_094 = data_d1[471:464];
        7'd60: vec_data_094 = data_d1[479:472];
        7'd61: vec_data_094 = data_d1[487:480];
        7'd62: vec_data_094 = data_d1[495:488];
        7'd63: vec_data_094 = data_d1[503:496];
        7'd64: vec_data_094 = data_d1[511:504];
        7'd65: vec_data_094 = data_d1[519:512];
        7'd66: vec_data_094 = data_d1[527:520];
        7'd67: vec_data_094 = data_d1[535:528];
        7'd68: vec_data_094 = data_d1[543:536];
        7'd69: vec_data_094 = data_d1[551:544];
        7'd70: vec_data_094 = data_d1[559:552];
        7'd71: vec_data_094 = data_d1[567:560];
        7'd72: vec_data_094 = data_d1[575:568];
        7'd73: vec_data_094 = data_d1[583:576];
        7'd74: vec_data_094 = data_d1[591:584];
        7'd75: vec_data_094 = data_d1[599:592];
        7'd76: vec_data_094 = data_d1[607:600];
        7'd77: vec_data_094 = data_d1[615:608];
        7'd78: vec_data_094 = data_d1[623:616];
        7'd79: vec_data_094 = data_d1[631:624];
        7'd80: vec_data_094 = data_d1[639:632];
        7'd81: vec_data_094 = data_d1[647:640];
        7'd82: vec_data_094 = data_d1[655:648];
        7'd83: vec_data_094 = data_d1[663:656];
        7'd84: vec_data_094 = data_d1[671:664];
        7'd85: vec_data_094 = data_d1[679:672];
        7'd86: vec_data_094 = data_d1[687:680];
        7'd87: vec_data_094 = data_d1[695:688];
        7'd88: vec_data_094 = data_d1[703:696];
        7'd89: vec_data_094 = data_d1[711:704];
        7'd90: vec_data_094 = data_d1[719:712];
        7'd91: vec_data_094 = data_d1[727:720];
        7'd92: vec_data_094 = data_d1[735:728];
        7'd93: vec_data_094 = data_d1[743:736];
        7'd94: vec_data_094 = data_d1[751:744];
        7'd95: vec_data_094 = data_d1[759:752];
    endcase
end

always @(
  vec_sum_095_d1
  or data_d1
  ) begin
    vec_data_095 = 8'b0;
    case(vec_sum_095_d1)
        7'd1: vec_data_095 = data_d1[7:0];
        7'd2: vec_data_095 = data_d1[15:8];
        7'd3: vec_data_095 = data_d1[23:16];
        7'd4: vec_data_095 = data_d1[31:24];
        7'd5: vec_data_095 = data_d1[39:32];
        7'd6: vec_data_095 = data_d1[47:40];
        7'd7: vec_data_095 = data_d1[55:48];
        7'd8: vec_data_095 = data_d1[63:56];
        7'd9: vec_data_095 = data_d1[71:64];
        7'd10: vec_data_095 = data_d1[79:72];
        7'd11: vec_data_095 = data_d1[87:80];
        7'd12: vec_data_095 = data_d1[95:88];
        7'd13: vec_data_095 = data_d1[103:96];
        7'd14: vec_data_095 = data_d1[111:104];
        7'd15: vec_data_095 = data_d1[119:112];
        7'd16: vec_data_095 = data_d1[127:120];
        7'd17: vec_data_095 = data_d1[135:128];
        7'd18: vec_data_095 = data_d1[143:136];
        7'd19: vec_data_095 = data_d1[151:144];
        7'd20: vec_data_095 = data_d1[159:152];
        7'd21: vec_data_095 = data_d1[167:160];
        7'd22: vec_data_095 = data_d1[175:168];
        7'd23: vec_data_095 = data_d1[183:176];
        7'd24: vec_data_095 = data_d1[191:184];
        7'd25: vec_data_095 = data_d1[199:192];
        7'd26: vec_data_095 = data_d1[207:200];
        7'd27: vec_data_095 = data_d1[215:208];
        7'd28: vec_data_095 = data_d1[223:216];
        7'd29: vec_data_095 = data_d1[231:224];
        7'd30: vec_data_095 = data_d1[239:232];
        7'd31: vec_data_095 = data_d1[247:240];
        7'd32: vec_data_095 = data_d1[255:248];
        7'd33: vec_data_095 = data_d1[263:256];
        7'd34: vec_data_095 = data_d1[271:264];
        7'd35: vec_data_095 = data_d1[279:272];
        7'd36: vec_data_095 = data_d1[287:280];
        7'd37: vec_data_095 = data_d1[295:288];
        7'd38: vec_data_095 = data_d1[303:296];
        7'd39: vec_data_095 = data_d1[311:304];
        7'd40: vec_data_095 = data_d1[319:312];
        7'd41: vec_data_095 = data_d1[327:320];
        7'd42: vec_data_095 = data_d1[335:328];
        7'd43: vec_data_095 = data_d1[343:336];
        7'd44: vec_data_095 = data_d1[351:344];
        7'd45: vec_data_095 = data_d1[359:352];
        7'd46: vec_data_095 = data_d1[367:360];
        7'd47: vec_data_095 = data_d1[375:368];
        7'd48: vec_data_095 = data_d1[383:376];
        7'd49: vec_data_095 = data_d1[391:384];
        7'd50: vec_data_095 = data_d1[399:392];
        7'd51: vec_data_095 = data_d1[407:400];
        7'd52: vec_data_095 = data_d1[415:408];
        7'd53: vec_data_095 = data_d1[423:416];
        7'd54: vec_data_095 = data_d1[431:424];
        7'd55: vec_data_095 = data_d1[439:432];
        7'd56: vec_data_095 = data_d1[447:440];
        7'd57: vec_data_095 = data_d1[455:448];
        7'd58: vec_data_095 = data_d1[463:456];
        7'd59: vec_data_095 = data_d1[471:464];
        7'd60: vec_data_095 = data_d1[479:472];
        7'd61: vec_data_095 = data_d1[487:480];
        7'd62: vec_data_095 = data_d1[495:488];
        7'd63: vec_data_095 = data_d1[503:496];
        7'd64: vec_data_095 = data_d1[511:504];
        7'd65: vec_data_095 = data_d1[519:512];
        7'd66: vec_data_095 = data_d1[527:520];
        7'd67: vec_data_095 = data_d1[535:528];
        7'd68: vec_data_095 = data_d1[543:536];
        7'd69: vec_data_095 = data_d1[551:544];
        7'd70: vec_data_095 = data_d1[559:552];
        7'd71: vec_data_095 = data_d1[567:560];
        7'd72: vec_data_095 = data_d1[575:568];
        7'd73: vec_data_095 = data_d1[583:576];
        7'd74: vec_data_095 = data_d1[591:584];
        7'd75: vec_data_095 = data_d1[599:592];
        7'd76: vec_data_095 = data_d1[607:600];
        7'd77: vec_data_095 = data_d1[615:608];
        7'd78: vec_data_095 = data_d1[623:616];
        7'd79: vec_data_095 = data_d1[631:624];
        7'd80: vec_data_095 = data_d1[639:632];
        7'd81: vec_data_095 = data_d1[647:640];
        7'd82: vec_data_095 = data_d1[655:648];
        7'd83: vec_data_095 = data_d1[663:656];
        7'd84: vec_data_095 = data_d1[671:664];
        7'd85: vec_data_095 = data_d1[679:672];
        7'd86: vec_data_095 = data_d1[687:680];
        7'd87: vec_data_095 = data_d1[695:688];
        7'd88: vec_data_095 = data_d1[703:696];
        7'd89: vec_data_095 = data_d1[711:704];
        7'd90: vec_data_095 = data_d1[719:712];
        7'd91: vec_data_095 = data_d1[727:720];
        7'd92: vec_data_095 = data_d1[735:728];
        7'd93: vec_data_095 = data_d1[743:736];
        7'd94: vec_data_095 = data_d1[751:744];
        7'd95: vec_data_095 = data_d1[759:752];
        7'd96: vec_data_095 = data_d1[767:760];
    endcase
end

always @(
  vec_sum_096_d1
  or data_d1
  ) begin
    vec_data_096 = 8'b0;
    case(vec_sum_096_d1)
        7'd1: vec_data_096 = data_d1[7:0];
        7'd2: vec_data_096 = data_d1[15:8];
        7'd3: vec_data_096 = data_d1[23:16];
        7'd4: vec_data_096 = data_d1[31:24];
        7'd5: vec_data_096 = data_d1[39:32];
        7'd6: vec_data_096 = data_d1[47:40];
        7'd7: vec_data_096 = data_d1[55:48];
        7'd8: vec_data_096 = data_d1[63:56];
        7'd9: vec_data_096 = data_d1[71:64];
        7'd10: vec_data_096 = data_d1[79:72];
        7'd11: vec_data_096 = data_d1[87:80];
        7'd12: vec_data_096 = data_d1[95:88];
        7'd13: vec_data_096 = data_d1[103:96];
        7'd14: vec_data_096 = data_d1[111:104];
        7'd15: vec_data_096 = data_d1[119:112];
        7'd16: vec_data_096 = data_d1[127:120];
        7'd17: vec_data_096 = data_d1[135:128];
        7'd18: vec_data_096 = data_d1[143:136];
        7'd19: vec_data_096 = data_d1[151:144];
        7'd20: vec_data_096 = data_d1[159:152];
        7'd21: vec_data_096 = data_d1[167:160];
        7'd22: vec_data_096 = data_d1[175:168];
        7'd23: vec_data_096 = data_d1[183:176];
        7'd24: vec_data_096 = data_d1[191:184];
        7'd25: vec_data_096 = data_d1[199:192];
        7'd26: vec_data_096 = data_d1[207:200];
        7'd27: vec_data_096 = data_d1[215:208];
        7'd28: vec_data_096 = data_d1[223:216];
        7'd29: vec_data_096 = data_d1[231:224];
        7'd30: vec_data_096 = data_d1[239:232];
        7'd31: vec_data_096 = data_d1[247:240];
        7'd32: vec_data_096 = data_d1[255:248];
        7'd33: vec_data_096 = data_d1[263:256];
        7'd34: vec_data_096 = data_d1[271:264];
        7'd35: vec_data_096 = data_d1[279:272];
        7'd36: vec_data_096 = data_d1[287:280];
        7'd37: vec_data_096 = data_d1[295:288];
        7'd38: vec_data_096 = data_d1[303:296];
        7'd39: vec_data_096 = data_d1[311:304];
        7'd40: vec_data_096 = data_d1[319:312];
        7'd41: vec_data_096 = data_d1[327:320];
        7'd42: vec_data_096 = data_d1[335:328];
        7'd43: vec_data_096 = data_d1[343:336];
        7'd44: vec_data_096 = data_d1[351:344];
        7'd45: vec_data_096 = data_d1[359:352];
        7'd46: vec_data_096 = data_d1[367:360];
        7'd47: vec_data_096 = data_d1[375:368];
        7'd48: vec_data_096 = data_d1[383:376];
        7'd49: vec_data_096 = data_d1[391:384];
        7'd50: vec_data_096 = data_d1[399:392];
        7'd51: vec_data_096 = data_d1[407:400];
        7'd52: vec_data_096 = data_d1[415:408];
        7'd53: vec_data_096 = data_d1[423:416];
        7'd54: vec_data_096 = data_d1[431:424];
        7'd55: vec_data_096 = data_d1[439:432];
        7'd56: vec_data_096 = data_d1[447:440];
        7'd57: vec_data_096 = data_d1[455:448];
        7'd58: vec_data_096 = data_d1[463:456];
        7'd59: vec_data_096 = data_d1[471:464];
        7'd60: vec_data_096 = data_d1[479:472];
        7'd61: vec_data_096 = data_d1[487:480];
        7'd62: vec_data_096 = data_d1[495:488];
        7'd63: vec_data_096 = data_d1[503:496];
        7'd64: vec_data_096 = data_d1[511:504];
        7'd65: vec_data_096 = data_d1[519:512];
        7'd66: vec_data_096 = data_d1[527:520];
        7'd67: vec_data_096 = data_d1[535:528];
        7'd68: vec_data_096 = data_d1[543:536];
        7'd69: vec_data_096 = data_d1[551:544];
        7'd70: vec_data_096 = data_d1[559:552];
        7'd71: vec_data_096 = data_d1[567:560];
        7'd72: vec_data_096 = data_d1[575:568];
        7'd73: vec_data_096 = data_d1[583:576];
        7'd74: vec_data_096 = data_d1[591:584];
        7'd75: vec_data_096 = data_d1[599:592];
        7'd76: vec_data_096 = data_d1[607:600];
        7'd77: vec_data_096 = data_d1[615:608];
        7'd78: vec_data_096 = data_d1[623:616];
        7'd79: vec_data_096 = data_d1[631:624];
        7'd80: vec_data_096 = data_d1[639:632];
        7'd81: vec_data_096 = data_d1[647:640];
        7'd82: vec_data_096 = data_d1[655:648];
        7'd83: vec_data_096 = data_d1[663:656];
        7'd84: vec_data_096 = data_d1[671:664];
        7'd85: vec_data_096 = data_d1[679:672];
        7'd86: vec_data_096 = data_d1[687:680];
        7'd87: vec_data_096 = data_d1[695:688];
        7'd88: vec_data_096 = data_d1[703:696];
        7'd89: vec_data_096 = data_d1[711:704];
        7'd90: vec_data_096 = data_d1[719:712];
        7'd91: vec_data_096 = data_d1[727:720];
        7'd92: vec_data_096 = data_d1[735:728];
        7'd93: vec_data_096 = data_d1[743:736];
        7'd94: vec_data_096 = data_d1[751:744];
        7'd95: vec_data_096 = data_d1[759:752];
        7'd96: vec_data_096 = data_d1[767:760];
        7'd97: vec_data_096 = data_d1[775:768];
    endcase
end

always @(
  vec_sum_097_d1
  or data_d1
  ) begin
    vec_data_097 = 8'b0;
    case(vec_sum_097_d1)
        7'd1: vec_data_097 = data_d1[7:0];
        7'd2: vec_data_097 = data_d1[15:8];
        7'd3: vec_data_097 = data_d1[23:16];
        7'd4: vec_data_097 = data_d1[31:24];
        7'd5: vec_data_097 = data_d1[39:32];
        7'd6: vec_data_097 = data_d1[47:40];
        7'd7: vec_data_097 = data_d1[55:48];
        7'd8: vec_data_097 = data_d1[63:56];
        7'd9: vec_data_097 = data_d1[71:64];
        7'd10: vec_data_097 = data_d1[79:72];
        7'd11: vec_data_097 = data_d1[87:80];
        7'd12: vec_data_097 = data_d1[95:88];
        7'd13: vec_data_097 = data_d1[103:96];
        7'd14: vec_data_097 = data_d1[111:104];
        7'd15: vec_data_097 = data_d1[119:112];
        7'd16: vec_data_097 = data_d1[127:120];
        7'd17: vec_data_097 = data_d1[135:128];
        7'd18: vec_data_097 = data_d1[143:136];
        7'd19: vec_data_097 = data_d1[151:144];
        7'd20: vec_data_097 = data_d1[159:152];
        7'd21: vec_data_097 = data_d1[167:160];
        7'd22: vec_data_097 = data_d1[175:168];
        7'd23: vec_data_097 = data_d1[183:176];
        7'd24: vec_data_097 = data_d1[191:184];
        7'd25: vec_data_097 = data_d1[199:192];
        7'd26: vec_data_097 = data_d1[207:200];
        7'd27: vec_data_097 = data_d1[215:208];
        7'd28: vec_data_097 = data_d1[223:216];
        7'd29: vec_data_097 = data_d1[231:224];
        7'd30: vec_data_097 = data_d1[239:232];
        7'd31: vec_data_097 = data_d1[247:240];
        7'd32: vec_data_097 = data_d1[255:248];
        7'd33: vec_data_097 = data_d1[263:256];
        7'd34: vec_data_097 = data_d1[271:264];
        7'd35: vec_data_097 = data_d1[279:272];
        7'd36: vec_data_097 = data_d1[287:280];
        7'd37: vec_data_097 = data_d1[295:288];
        7'd38: vec_data_097 = data_d1[303:296];
        7'd39: vec_data_097 = data_d1[311:304];
        7'd40: vec_data_097 = data_d1[319:312];
        7'd41: vec_data_097 = data_d1[327:320];
        7'd42: vec_data_097 = data_d1[335:328];
        7'd43: vec_data_097 = data_d1[343:336];
        7'd44: vec_data_097 = data_d1[351:344];
        7'd45: vec_data_097 = data_d1[359:352];
        7'd46: vec_data_097 = data_d1[367:360];
        7'd47: vec_data_097 = data_d1[375:368];
        7'd48: vec_data_097 = data_d1[383:376];
        7'd49: vec_data_097 = data_d1[391:384];
        7'd50: vec_data_097 = data_d1[399:392];
        7'd51: vec_data_097 = data_d1[407:400];
        7'd52: vec_data_097 = data_d1[415:408];
        7'd53: vec_data_097 = data_d1[423:416];
        7'd54: vec_data_097 = data_d1[431:424];
        7'd55: vec_data_097 = data_d1[439:432];
        7'd56: vec_data_097 = data_d1[447:440];
        7'd57: vec_data_097 = data_d1[455:448];
        7'd58: vec_data_097 = data_d1[463:456];
        7'd59: vec_data_097 = data_d1[471:464];
        7'd60: vec_data_097 = data_d1[479:472];
        7'd61: vec_data_097 = data_d1[487:480];
        7'd62: vec_data_097 = data_d1[495:488];
        7'd63: vec_data_097 = data_d1[503:496];
        7'd64: vec_data_097 = data_d1[511:504];
        7'd65: vec_data_097 = data_d1[519:512];
        7'd66: vec_data_097 = data_d1[527:520];
        7'd67: vec_data_097 = data_d1[535:528];
        7'd68: vec_data_097 = data_d1[543:536];
        7'd69: vec_data_097 = data_d1[551:544];
        7'd70: vec_data_097 = data_d1[559:552];
        7'd71: vec_data_097 = data_d1[567:560];
        7'd72: vec_data_097 = data_d1[575:568];
        7'd73: vec_data_097 = data_d1[583:576];
        7'd74: vec_data_097 = data_d1[591:584];
        7'd75: vec_data_097 = data_d1[599:592];
        7'd76: vec_data_097 = data_d1[607:600];
        7'd77: vec_data_097 = data_d1[615:608];
        7'd78: vec_data_097 = data_d1[623:616];
        7'd79: vec_data_097 = data_d1[631:624];
        7'd80: vec_data_097 = data_d1[639:632];
        7'd81: vec_data_097 = data_d1[647:640];
        7'd82: vec_data_097 = data_d1[655:648];
        7'd83: vec_data_097 = data_d1[663:656];
        7'd84: vec_data_097 = data_d1[671:664];
        7'd85: vec_data_097 = data_d1[679:672];
        7'd86: vec_data_097 = data_d1[687:680];
        7'd87: vec_data_097 = data_d1[695:688];
        7'd88: vec_data_097 = data_d1[703:696];
        7'd89: vec_data_097 = data_d1[711:704];
        7'd90: vec_data_097 = data_d1[719:712];
        7'd91: vec_data_097 = data_d1[727:720];
        7'd92: vec_data_097 = data_d1[735:728];
        7'd93: vec_data_097 = data_d1[743:736];
        7'd94: vec_data_097 = data_d1[751:744];
        7'd95: vec_data_097 = data_d1[759:752];
        7'd96: vec_data_097 = data_d1[767:760];
        7'd97: vec_data_097 = data_d1[775:768];
        7'd98: vec_data_097 = data_d1[783:776];
    endcase
end

always @(
  vec_sum_098_d1
  or data_d1
  ) begin
    vec_data_098 = 8'b0;
    case(vec_sum_098_d1)
        7'd1: vec_data_098 = data_d1[7:0];
        7'd2: vec_data_098 = data_d1[15:8];
        7'd3: vec_data_098 = data_d1[23:16];
        7'd4: vec_data_098 = data_d1[31:24];
        7'd5: vec_data_098 = data_d1[39:32];
        7'd6: vec_data_098 = data_d1[47:40];
        7'd7: vec_data_098 = data_d1[55:48];
        7'd8: vec_data_098 = data_d1[63:56];
        7'd9: vec_data_098 = data_d1[71:64];
        7'd10: vec_data_098 = data_d1[79:72];
        7'd11: vec_data_098 = data_d1[87:80];
        7'd12: vec_data_098 = data_d1[95:88];
        7'd13: vec_data_098 = data_d1[103:96];
        7'd14: vec_data_098 = data_d1[111:104];
        7'd15: vec_data_098 = data_d1[119:112];
        7'd16: vec_data_098 = data_d1[127:120];
        7'd17: vec_data_098 = data_d1[135:128];
        7'd18: vec_data_098 = data_d1[143:136];
        7'd19: vec_data_098 = data_d1[151:144];
        7'd20: vec_data_098 = data_d1[159:152];
        7'd21: vec_data_098 = data_d1[167:160];
        7'd22: vec_data_098 = data_d1[175:168];
        7'd23: vec_data_098 = data_d1[183:176];
        7'd24: vec_data_098 = data_d1[191:184];
        7'd25: vec_data_098 = data_d1[199:192];
        7'd26: vec_data_098 = data_d1[207:200];
        7'd27: vec_data_098 = data_d1[215:208];
        7'd28: vec_data_098 = data_d1[223:216];
        7'd29: vec_data_098 = data_d1[231:224];
        7'd30: vec_data_098 = data_d1[239:232];
        7'd31: vec_data_098 = data_d1[247:240];
        7'd32: vec_data_098 = data_d1[255:248];
        7'd33: vec_data_098 = data_d1[263:256];
        7'd34: vec_data_098 = data_d1[271:264];
        7'd35: vec_data_098 = data_d1[279:272];
        7'd36: vec_data_098 = data_d1[287:280];
        7'd37: vec_data_098 = data_d1[295:288];
        7'd38: vec_data_098 = data_d1[303:296];
        7'd39: vec_data_098 = data_d1[311:304];
        7'd40: vec_data_098 = data_d1[319:312];
        7'd41: vec_data_098 = data_d1[327:320];
        7'd42: vec_data_098 = data_d1[335:328];
        7'd43: vec_data_098 = data_d1[343:336];
        7'd44: vec_data_098 = data_d1[351:344];
        7'd45: vec_data_098 = data_d1[359:352];
        7'd46: vec_data_098 = data_d1[367:360];
        7'd47: vec_data_098 = data_d1[375:368];
        7'd48: vec_data_098 = data_d1[383:376];
        7'd49: vec_data_098 = data_d1[391:384];
        7'd50: vec_data_098 = data_d1[399:392];
        7'd51: vec_data_098 = data_d1[407:400];
        7'd52: vec_data_098 = data_d1[415:408];
        7'd53: vec_data_098 = data_d1[423:416];
        7'd54: vec_data_098 = data_d1[431:424];
        7'd55: vec_data_098 = data_d1[439:432];
        7'd56: vec_data_098 = data_d1[447:440];
        7'd57: vec_data_098 = data_d1[455:448];
        7'd58: vec_data_098 = data_d1[463:456];
        7'd59: vec_data_098 = data_d1[471:464];
        7'd60: vec_data_098 = data_d1[479:472];
        7'd61: vec_data_098 = data_d1[487:480];
        7'd62: vec_data_098 = data_d1[495:488];
        7'd63: vec_data_098 = data_d1[503:496];
        7'd64: vec_data_098 = data_d1[511:504];
        7'd65: vec_data_098 = data_d1[519:512];
        7'd66: vec_data_098 = data_d1[527:520];
        7'd67: vec_data_098 = data_d1[535:528];
        7'd68: vec_data_098 = data_d1[543:536];
        7'd69: vec_data_098 = data_d1[551:544];
        7'd70: vec_data_098 = data_d1[559:552];
        7'd71: vec_data_098 = data_d1[567:560];
        7'd72: vec_data_098 = data_d1[575:568];
        7'd73: vec_data_098 = data_d1[583:576];
        7'd74: vec_data_098 = data_d1[591:584];
        7'd75: vec_data_098 = data_d1[599:592];
        7'd76: vec_data_098 = data_d1[607:600];
        7'd77: vec_data_098 = data_d1[615:608];
        7'd78: vec_data_098 = data_d1[623:616];
        7'd79: vec_data_098 = data_d1[631:624];
        7'd80: vec_data_098 = data_d1[639:632];
        7'd81: vec_data_098 = data_d1[647:640];
        7'd82: vec_data_098 = data_d1[655:648];
        7'd83: vec_data_098 = data_d1[663:656];
        7'd84: vec_data_098 = data_d1[671:664];
        7'd85: vec_data_098 = data_d1[679:672];
        7'd86: vec_data_098 = data_d1[687:680];
        7'd87: vec_data_098 = data_d1[695:688];
        7'd88: vec_data_098 = data_d1[703:696];
        7'd89: vec_data_098 = data_d1[711:704];
        7'd90: vec_data_098 = data_d1[719:712];
        7'd91: vec_data_098 = data_d1[727:720];
        7'd92: vec_data_098 = data_d1[735:728];
        7'd93: vec_data_098 = data_d1[743:736];
        7'd94: vec_data_098 = data_d1[751:744];
        7'd95: vec_data_098 = data_d1[759:752];
        7'd96: vec_data_098 = data_d1[767:760];
        7'd97: vec_data_098 = data_d1[775:768];
        7'd98: vec_data_098 = data_d1[783:776];
        7'd99: vec_data_098 = data_d1[791:784];
    endcase
end

always @(
  vec_sum_099_d1
  or data_d1
  ) begin
    vec_data_099 = 8'b0;
    case(vec_sum_099_d1)
        7'd1: vec_data_099 = data_d1[7:0];
        7'd2: vec_data_099 = data_d1[15:8];
        7'd3: vec_data_099 = data_d1[23:16];
        7'd4: vec_data_099 = data_d1[31:24];
        7'd5: vec_data_099 = data_d1[39:32];
        7'd6: vec_data_099 = data_d1[47:40];
        7'd7: vec_data_099 = data_d1[55:48];
        7'd8: vec_data_099 = data_d1[63:56];
        7'd9: vec_data_099 = data_d1[71:64];
        7'd10: vec_data_099 = data_d1[79:72];
        7'd11: vec_data_099 = data_d1[87:80];
        7'd12: vec_data_099 = data_d1[95:88];
        7'd13: vec_data_099 = data_d1[103:96];
        7'd14: vec_data_099 = data_d1[111:104];
        7'd15: vec_data_099 = data_d1[119:112];
        7'd16: vec_data_099 = data_d1[127:120];
        7'd17: vec_data_099 = data_d1[135:128];
        7'd18: vec_data_099 = data_d1[143:136];
        7'd19: vec_data_099 = data_d1[151:144];
        7'd20: vec_data_099 = data_d1[159:152];
        7'd21: vec_data_099 = data_d1[167:160];
        7'd22: vec_data_099 = data_d1[175:168];
        7'd23: vec_data_099 = data_d1[183:176];
        7'd24: vec_data_099 = data_d1[191:184];
        7'd25: vec_data_099 = data_d1[199:192];
        7'd26: vec_data_099 = data_d1[207:200];
        7'd27: vec_data_099 = data_d1[215:208];
        7'd28: vec_data_099 = data_d1[223:216];
        7'd29: vec_data_099 = data_d1[231:224];
        7'd30: vec_data_099 = data_d1[239:232];
        7'd31: vec_data_099 = data_d1[247:240];
        7'd32: vec_data_099 = data_d1[255:248];
        7'd33: vec_data_099 = data_d1[263:256];
        7'd34: vec_data_099 = data_d1[271:264];
        7'd35: vec_data_099 = data_d1[279:272];
        7'd36: vec_data_099 = data_d1[287:280];
        7'd37: vec_data_099 = data_d1[295:288];
        7'd38: vec_data_099 = data_d1[303:296];
        7'd39: vec_data_099 = data_d1[311:304];
        7'd40: vec_data_099 = data_d1[319:312];
        7'd41: vec_data_099 = data_d1[327:320];
        7'd42: vec_data_099 = data_d1[335:328];
        7'd43: vec_data_099 = data_d1[343:336];
        7'd44: vec_data_099 = data_d1[351:344];
        7'd45: vec_data_099 = data_d1[359:352];
        7'd46: vec_data_099 = data_d1[367:360];
        7'd47: vec_data_099 = data_d1[375:368];
        7'd48: vec_data_099 = data_d1[383:376];
        7'd49: vec_data_099 = data_d1[391:384];
        7'd50: vec_data_099 = data_d1[399:392];
        7'd51: vec_data_099 = data_d1[407:400];
        7'd52: vec_data_099 = data_d1[415:408];
        7'd53: vec_data_099 = data_d1[423:416];
        7'd54: vec_data_099 = data_d1[431:424];
        7'd55: vec_data_099 = data_d1[439:432];
        7'd56: vec_data_099 = data_d1[447:440];
        7'd57: vec_data_099 = data_d1[455:448];
        7'd58: vec_data_099 = data_d1[463:456];
        7'd59: vec_data_099 = data_d1[471:464];
        7'd60: vec_data_099 = data_d1[479:472];
        7'd61: vec_data_099 = data_d1[487:480];
        7'd62: vec_data_099 = data_d1[495:488];
        7'd63: vec_data_099 = data_d1[503:496];
        7'd64: vec_data_099 = data_d1[511:504];
        7'd65: vec_data_099 = data_d1[519:512];
        7'd66: vec_data_099 = data_d1[527:520];
        7'd67: vec_data_099 = data_d1[535:528];
        7'd68: vec_data_099 = data_d1[543:536];
        7'd69: vec_data_099 = data_d1[551:544];
        7'd70: vec_data_099 = data_d1[559:552];
        7'd71: vec_data_099 = data_d1[567:560];
        7'd72: vec_data_099 = data_d1[575:568];
        7'd73: vec_data_099 = data_d1[583:576];
        7'd74: vec_data_099 = data_d1[591:584];
        7'd75: vec_data_099 = data_d1[599:592];
        7'd76: vec_data_099 = data_d1[607:600];
        7'd77: vec_data_099 = data_d1[615:608];
        7'd78: vec_data_099 = data_d1[623:616];
        7'd79: vec_data_099 = data_d1[631:624];
        7'd80: vec_data_099 = data_d1[639:632];
        7'd81: vec_data_099 = data_d1[647:640];
        7'd82: vec_data_099 = data_d1[655:648];
        7'd83: vec_data_099 = data_d1[663:656];
        7'd84: vec_data_099 = data_d1[671:664];
        7'd85: vec_data_099 = data_d1[679:672];
        7'd86: vec_data_099 = data_d1[687:680];
        7'd87: vec_data_099 = data_d1[695:688];
        7'd88: vec_data_099 = data_d1[703:696];
        7'd89: vec_data_099 = data_d1[711:704];
        7'd90: vec_data_099 = data_d1[719:712];
        7'd91: vec_data_099 = data_d1[727:720];
        7'd92: vec_data_099 = data_d1[735:728];
        7'd93: vec_data_099 = data_d1[743:736];
        7'd94: vec_data_099 = data_d1[751:744];
        7'd95: vec_data_099 = data_d1[759:752];
        7'd96: vec_data_099 = data_d1[767:760];
        7'd97: vec_data_099 = data_d1[775:768];
        7'd98: vec_data_099 = data_d1[783:776];
        7'd99: vec_data_099 = data_d1[791:784];
        7'd100: vec_data_099 = data_d1[799:792];
    endcase
end

always @(
  vec_sum_100_d1
  or data_d1
  ) begin
    vec_data_100 = 8'b0;
    case(vec_sum_100_d1)
        7'd1: vec_data_100 = data_d1[7:0];
        7'd2: vec_data_100 = data_d1[15:8];
        7'd3: vec_data_100 = data_d1[23:16];
        7'd4: vec_data_100 = data_d1[31:24];
        7'd5: vec_data_100 = data_d1[39:32];
        7'd6: vec_data_100 = data_d1[47:40];
        7'd7: vec_data_100 = data_d1[55:48];
        7'd8: vec_data_100 = data_d1[63:56];
        7'd9: vec_data_100 = data_d1[71:64];
        7'd10: vec_data_100 = data_d1[79:72];
        7'd11: vec_data_100 = data_d1[87:80];
        7'd12: vec_data_100 = data_d1[95:88];
        7'd13: vec_data_100 = data_d1[103:96];
        7'd14: vec_data_100 = data_d1[111:104];
        7'd15: vec_data_100 = data_d1[119:112];
        7'd16: vec_data_100 = data_d1[127:120];
        7'd17: vec_data_100 = data_d1[135:128];
        7'd18: vec_data_100 = data_d1[143:136];
        7'd19: vec_data_100 = data_d1[151:144];
        7'd20: vec_data_100 = data_d1[159:152];
        7'd21: vec_data_100 = data_d1[167:160];
        7'd22: vec_data_100 = data_d1[175:168];
        7'd23: vec_data_100 = data_d1[183:176];
        7'd24: vec_data_100 = data_d1[191:184];
        7'd25: vec_data_100 = data_d1[199:192];
        7'd26: vec_data_100 = data_d1[207:200];
        7'd27: vec_data_100 = data_d1[215:208];
        7'd28: vec_data_100 = data_d1[223:216];
        7'd29: vec_data_100 = data_d1[231:224];
        7'd30: vec_data_100 = data_d1[239:232];
        7'd31: vec_data_100 = data_d1[247:240];
        7'd32: vec_data_100 = data_d1[255:248];
        7'd33: vec_data_100 = data_d1[263:256];
        7'd34: vec_data_100 = data_d1[271:264];
        7'd35: vec_data_100 = data_d1[279:272];
        7'd36: vec_data_100 = data_d1[287:280];
        7'd37: vec_data_100 = data_d1[295:288];
        7'd38: vec_data_100 = data_d1[303:296];
        7'd39: vec_data_100 = data_d1[311:304];
        7'd40: vec_data_100 = data_d1[319:312];
        7'd41: vec_data_100 = data_d1[327:320];
        7'd42: vec_data_100 = data_d1[335:328];
        7'd43: vec_data_100 = data_d1[343:336];
        7'd44: vec_data_100 = data_d1[351:344];
        7'd45: vec_data_100 = data_d1[359:352];
        7'd46: vec_data_100 = data_d1[367:360];
        7'd47: vec_data_100 = data_d1[375:368];
        7'd48: vec_data_100 = data_d1[383:376];
        7'd49: vec_data_100 = data_d1[391:384];
        7'd50: vec_data_100 = data_d1[399:392];
        7'd51: vec_data_100 = data_d1[407:400];
        7'd52: vec_data_100 = data_d1[415:408];
        7'd53: vec_data_100 = data_d1[423:416];
        7'd54: vec_data_100 = data_d1[431:424];
        7'd55: vec_data_100 = data_d1[439:432];
        7'd56: vec_data_100 = data_d1[447:440];
        7'd57: vec_data_100 = data_d1[455:448];
        7'd58: vec_data_100 = data_d1[463:456];
        7'd59: vec_data_100 = data_d1[471:464];
        7'd60: vec_data_100 = data_d1[479:472];
        7'd61: vec_data_100 = data_d1[487:480];
        7'd62: vec_data_100 = data_d1[495:488];
        7'd63: vec_data_100 = data_d1[503:496];
        7'd64: vec_data_100 = data_d1[511:504];
        7'd65: vec_data_100 = data_d1[519:512];
        7'd66: vec_data_100 = data_d1[527:520];
        7'd67: vec_data_100 = data_d1[535:528];
        7'd68: vec_data_100 = data_d1[543:536];
        7'd69: vec_data_100 = data_d1[551:544];
        7'd70: vec_data_100 = data_d1[559:552];
        7'd71: vec_data_100 = data_d1[567:560];
        7'd72: vec_data_100 = data_d1[575:568];
        7'd73: vec_data_100 = data_d1[583:576];
        7'd74: vec_data_100 = data_d1[591:584];
        7'd75: vec_data_100 = data_d1[599:592];
        7'd76: vec_data_100 = data_d1[607:600];
        7'd77: vec_data_100 = data_d1[615:608];
        7'd78: vec_data_100 = data_d1[623:616];
        7'd79: vec_data_100 = data_d1[631:624];
        7'd80: vec_data_100 = data_d1[639:632];
        7'd81: vec_data_100 = data_d1[647:640];
        7'd82: vec_data_100 = data_d1[655:648];
        7'd83: vec_data_100 = data_d1[663:656];
        7'd84: vec_data_100 = data_d1[671:664];
        7'd85: vec_data_100 = data_d1[679:672];
        7'd86: vec_data_100 = data_d1[687:680];
        7'd87: vec_data_100 = data_d1[695:688];
        7'd88: vec_data_100 = data_d1[703:696];
        7'd89: vec_data_100 = data_d1[711:704];
        7'd90: vec_data_100 = data_d1[719:712];
        7'd91: vec_data_100 = data_d1[727:720];
        7'd92: vec_data_100 = data_d1[735:728];
        7'd93: vec_data_100 = data_d1[743:736];
        7'd94: vec_data_100 = data_d1[751:744];
        7'd95: vec_data_100 = data_d1[759:752];
        7'd96: vec_data_100 = data_d1[767:760];
        7'd97: vec_data_100 = data_d1[775:768];
        7'd98: vec_data_100 = data_d1[783:776];
        7'd99: vec_data_100 = data_d1[791:784];
        7'd100: vec_data_100 = data_d1[799:792];
        7'd101: vec_data_100 = data_d1[807:800];
    endcase
end

always @(
  vec_sum_101_d1
  or data_d1
  ) begin
    vec_data_101 = 8'b0;
    case(vec_sum_101_d1)
        7'd1: vec_data_101 = data_d1[7:0];
        7'd2: vec_data_101 = data_d1[15:8];
        7'd3: vec_data_101 = data_d1[23:16];
        7'd4: vec_data_101 = data_d1[31:24];
        7'd5: vec_data_101 = data_d1[39:32];
        7'd6: vec_data_101 = data_d1[47:40];
        7'd7: vec_data_101 = data_d1[55:48];
        7'd8: vec_data_101 = data_d1[63:56];
        7'd9: vec_data_101 = data_d1[71:64];
        7'd10: vec_data_101 = data_d1[79:72];
        7'd11: vec_data_101 = data_d1[87:80];
        7'd12: vec_data_101 = data_d1[95:88];
        7'd13: vec_data_101 = data_d1[103:96];
        7'd14: vec_data_101 = data_d1[111:104];
        7'd15: vec_data_101 = data_d1[119:112];
        7'd16: vec_data_101 = data_d1[127:120];
        7'd17: vec_data_101 = data_d1[135:128];
        7'd18: vec_data_101 = data_d1[143:136];
        7'd19: vec_data_101 = data_d1[151:144];
        7'd20: vec_data_101 = data_d1[159:152];
        7'd21: vec_data_101 = data_d1[167:160];
        7'd22: vec_data_101 = data_d1[175:168];
        7'd23: vec_data_101 = data_d1[183:176];
        7'd24: vec_data_101 = data_d1[191:184];
        7'd25: vec_data_101 = data_d1[199:192];
        7'd26: vec_data_101 = data_d1[207:200];
        7'd27: vec_data_101 = data_d1[215:208];
        7'd28: vec_data_101 = data_d1[223:216];
        7'd29: vec_data_101 = data_d1[231:224];
        7'd30: vec_data_101 = data_d1[239:232];
        7'd31: vec_data_101 = data_d1[247:240];
        7'd32: vec_data_101 = data_d1[255:248];
        7'd33: vec_data_101 = data_d1[263:256];
        7'd34: vec_data_101 = data_d1[271:264];
        7'd35: vec_data_101 = data_d1[279:272];
        7'd36: vec_data_101 = data_d1[287:280];
        7'd37: vec_data_101 = data_d1[295:288];
        7'd38: vec_data_101 = data_d1[303:296];
        7'd39: vec_data_101 = data_d1[311:304];
        7'd40: vec_data_101 = data_d1[319:312];
        7'd41: vec_data_101 = data_d1[327:320];
        7'd42: vec_data_101 = data_d1[335:328];
        7'd43: vec_data_101 = data_d1[343:336];
        7'd44: vec_data_101 = data_d1[351:344];
        7'd45: vec_data_101 = data_d1[359:352];
        7'd46: vec_data_101 = data_d1[367:360];
        7'd47: vec_data_101 = data_d1[375:368];
        7'd48: vec_data_101 = data_d1[383:376];
        7'd49: vec_data_101 = data_d1[391:384];
        7'd50: vec_data_101 = data_d1[399:392];
        7'd51: vec_data_101 = data_d1[407:400];
        7'd52: vec_data_101 = data_d1[415:408];
        7'd53: vec_data_101 = data_d1[423:416];
        7'd54: vec_data_101 = data_d1[431:424];
        7'd55: vec_data_101 = data_d1[439:432];
        7'd56: vec_data_101 = data_d1[447:440];
        7'd57: vec_data_101 = data_d1[455:448];
        7'd58: vec_data_101 = data_d1[463:456];
        7'd59: vec_data_101 = data_d1[471:464];
        7'd60: vec_data_101 = data_d1[479:472];
        7'd61: vec_data_101 = data_d1[487:480];
        7'd62: vec_data_101 = data_d1[495:488];
        7'd63: vec_data_101 = data_d1[503:496];
        7'd64: vec_data_101 = data_d1[511:504];
        7'd65: vec_data_101 = data_d1[519:512];
        7'd66: vec_data_101 = data_d1[527:520];
        7'd67: vec_data_101 = data_d1[535:528];
        7'd68: vec_data_101 = data_d1[543:536];
        7'd69: vec_data_101 = data_d1[551:544];
        7'd70: vec_data_101 = data_d1[559:552];
        7'd71: vec_data_101 = data_d1[567:560];
        7'd72: vec_data_101 = data_d1[575:568];
        7'd73: vec_data_101 = data_d1[583:576];
        7'd74: vec_data_101 = data_d1[591:584];
        7'd75: vec_data_101 = data_d1[599:592];
        7'd76: vec_data_101 = data_d1[607:600];
        7'd77: vec_data_101 = data_d1[615:608];
        7'd78: vec_data_101 = data_d1[623:616];
        7'd79: vec_data_101 = data_d1[631:624];
        7'd80: vec_data_101 = data_d1[639:632];
        7'd81: vec_data_101 = data_d1[647:640];
        7'd82: vec_data_101 = data_d1[655:648];
        7'd83: vec_data_101 = data_d1[663:656];
        7'd84: vec_data_101 = data_d1[671:664];
        7'd85: vec_data_101 = data_d1[679:672];
        7'd86: vec_data_101 = data_d1[687:680];
        7'd87: vec_data_101 = data_d1[695:688];
        7'd88: vec_data_101 = data_d1[703:696];
        7'd89: vec_data_101 = data_d1[711:704];
        7'd90: vec_data_101 = data_d1[719:712];
        7'd91: vec_data_101 = data_d1[727:720];
        7'd92: vec_data_101 = data_d1[735:728];
        7'd93: vec_data_101 = data_d1[743:736];
        7'd94: vec_data_101 = data_d1[751:744];
        7'd95: vec_data_101 = data_d1[759:752];
        7'd96: vec_data_101 = data_d1[767:760];
        7'd97: vec_data_101 = data_d1[775:768];
        7'd98: vec_data_101 = data_d1[783:776];
        7'd99: vec_data_101 = data_d1[791:784];
        7'd100: vec_data_101 = data_d1[799:792];
        7'd101: vec_data_101 = data_d1[807:800];
        7'd102: vec_data_101 = data_d1[815:808];
    endcase
end

always @(
  vec_sum_102_d1
  or data_d1
  ) begin
    vec_data_102 = 8'b0;
    case(vec_sum_102_d1)
        7'd1: vec_data_102 = data_d1[7:0];
        7'd2: vec_data_102 = data_d1[15:8];
        7'd3: vec_data_102 = data_d1[23:16];
        7'd4: vec_data_102 = data_d1[31:24];
        7'd5: vec_data_102 = data_d1[39:32];
        7'd6: vec_data_102 = data_d1[47:40];
        7'd7: vec_data_102 = data_d1[55:48];
        7'd8: vec_data_102 = data_d1[63:56];
        7'd9: vec_data_102 = data_d1[71:64];
        7'd10: vec_data_102 = data_d1[79:72];
        7'd11: vec_data_102 = data_d1[87:80];
        7'd12: vec_data_102 = data_d1[95:88];
        7'd13: vec_data_102 = data_d1[103:96];
        7'd14: vec_data_102 = data_d1[111:104];
        7'd15: vec_data_102 = data_d1[119:112];
        7'd16: vec_data_102 = data_d1[127:120];
        7'd17: vec_data_102 = data_d1[135:128];
        7'd18: vec_data_102 = data_d1[143:136];
        7'd19: vec_data_102 = data_d1[151:144];
        7'd20: vec_data_102 = data_d1[159:152];
        7'd21: vec_data_102 = data_d1[167:160];
        7'd22: vec_data_102 = data_d1[175:168];
        7'd23: vec_data_102 = data_d1[183:176];
        7'd24: vec_data_102 = data_d1[191:184];
        7'd25: vec_data_102 = data_d1[199:192];
        7'd26: vec_data_102 = data_d1[207:200];
        7'd27: vec_data_102 = data_d1[215:208];
        7'd28: vec_data_102 = data_d1[223:216];
        7'd29: vec_data_102 = data_d1[231:224];
        7'd30: vec_data_102 = data_d1[239:232];
        7'd31: vec_data_102 = data_d1[247:240];
        7'd32: vec_data_102 = data_d1[255:248];
        7'd33: vec_data_102 = data_d1[263:256];
        7'd34: vec_data_102 = data_d1[271:264];
        7'd35: vec_data_102 = data_d1[279:272];
        7'd36: vec_data_102 = data_d1[287:280];
        7'd37: vec_data_102 = data_d1[295:288];
        7'd38: vec_data_102 = data_d1[303:296];
        7'd39: vec_data_102 = data_d1[311:304];
        7'd40: vec_data_102 = data_d1[319:312];
        7'd41: vec_data_102 = data_d1[327:320];
        7'd42: vec_data_102 = data_d1[335:328];
        7'd43: vec_data_102 = data_d1[343:336];
        7'd44: vec_data_102 = data_d1[351:344];
        7'd45: vec_data_102 = data_d1[359:352];
        7'd46: vec_data_102 = data_d1[367:360];
        7'd47: vec_data_102 = data_d1[375:368];
        7'd48: vec_data_102 = data_d1[383:376];
        7'd49: vec_data_102 = data_d1[391:384];
        7'd50: vec_data_102 = data_d1[399:392];
        7'd51: vec_data_102 = data_d1[407:400];
        7'd52: vec_data_102 = data_d1[415:408];
        7'd53: vec_data_102 = data_d1[423:416];
        7'd54: vec_data_102 = data_d1[431:424];
        7'd55: vec_data_102 = data_d1[439:432];
        7'd56: vec_data_102 = data_d1[447:440];
        7'd57: vec_data_102 = data_d1[455:448];
        7'd58: vec_data_102 = data_d1[463:456];
        7'd59: vec_data_102 = data_d1[471:464];
        7'd60: vec_data_102 = data_d1[479:472];
        7'd61: vec_data_102 = data_d1[487:480];
        7'd62: vec_data_102 = data_d1[495:488];
        7'd63: vec_data_102 = data_d1[503:496];
        7'd64: vec_data_102 = data_d1[511:504];
        7'd65: vec_data_102 = data_d1[519:512];
        7'd66: vec_data_102 = data_d1[527:520];
        7'd67: vec_data_102 = data_d1[535:528];
        7'd68: vec_data_102 = data_d1[543:536];
        7'd69: vec_data_102 = data_d1[551:544];
        7'd70: vec_data_102 = data_d1[559:552];
        7'd71: vec_data_102 = data_d1[567:560];
        7'd72: vec_data_102 = data_d1[575:568];
        7'd73: vec_data_102 = data_d1[583:576];
        7'd74: vec_data_102 = data_d1[591:584];
        7'd75: vec_data_102 = data_d1[599:592];
        7'd76: vec_data_102 = data_d1[607:600];
        7'd77: vec_data_102 = data_d1[615:608];
        7'd78: vec_data_102 = data_d1[623:616];
        7'd79: vec_data_102 = data_d1[631:624];
        7'd80: vec_data_102 = data_d1[639:632];
        7'd81: vec_data_102 = data_d1[647:640];
        7'd82: vec_data_102 = data_d1[655:648];
        7'd83: vec_data_102 = data_d1[663:656];
        7'd84: vec_data_102 = data_d1[671:664];
        7'd85: vec_data_102 = data_d1[679:672];
        7'd86: vec_data_102 = data_d1[687:680];
        7'd87: vec_data_102 = data_d1[695:688];
        7'd88: vec_data_102 = data_d1[703:696];
        7'd89: vec_data_102 = data_d1[711:704];
        7'd90: vec_data_102 = data_d1[719:712];
        7'd91: vec_data_102 = data_d1[727:720];
        7'd92: vec_data_102 = data_d1[735:728];
        7'd93: vec_data_102 = data_d1[743:736];
        7'd94: vec_data_102 = data_d1[751:744];
        7'd95: vec_data_102 = data_d1[759:752];
        7'd96: vec_data_102 = data_d1[767:760];
        7'd97: vec_data_102 = data_d1[775:768];
        7'd98: vec_data_102 = data_d1[783:776];
        7'd99: vec_data_102 = data_d1[791:784];
        7'd100: vec_data_102 = data_d1[799:792];
        7'd101: vec_data_102 = data_d1[807:800];
        7'd102: vec_data_102 = data_d1[815:808];
        7'd103: vec_data_102 = data_d1[823:816];
    endcase
end

always @(
  vec_sum_103_d1
  or data_d1
  ) begin
    vec_data_103 = 8'b0;
    case(vec_sum_103_d1)
        7'd1: vec_data_103 = data_d1[7:0];
        7'd2: vec_data_103 = data_d1[15:8];
        7'd3: vec_data_103 = data_d1[23:16];
        7'd4: vec_data_103 = data_d1[31:24];
        7'd5: vec_data_103 = data_d1[39:32];
        7'd6: vec_data_103 = data_d1[47:40];
        7'd7: vec_data_103 = data_d1[55:48];
        7'd8: vec_data_103 = data_d1[63:56];
        7'd9: vec_data_103 = data_d1[71:64];
        7'd10: vec_data_103 = data_d1[79:72];
        7'd11: vec_data_103 = data_d1[87:80];
        7'd12: vec_data_103 = data_d1[95:88];
        7'd13: vec_data_103 = data_d1[103:96];
        7'd14: vec_data_103 = data_d1[111:104];
        7'd15: vec_data_103 = data_d1[119:112];
        7'd16: vec_data_103 = data_d1[127:120];
        7'd17: vec_data_103 = data_d1[135:128];
        7'd18: vec_data_103 = data_d1[143:136];
        7'd19: vec_data_103 = data_d1[151:144];
        7'd20: vec_data_103 = data_d1[159:152];
        7'd21: vec_data_103 = data_d1[167:160];
        7'd22: vec_data_103 = data_d1[175:168];
        7'd23: vec_data_103 = data_d1[183:176];
        7'd24: vec_data_103 = data_d1[191:184];
        7'd25: vec_data_103 = data_d1[199:192];
        7'd26: vec_data_103 = data_d1[207:200];
        7'd27: vec_data_103 = data_d1[215:208];
        7'd28: vec_data_103 = data_d1[223:216];
        7'd29: vec_data_103 = data_d1[231:224];
        7'd30: vec_data_103 = data_d1[239:232];
        7'd31: vec_data_103 = data_d1[247:240];
        7'd32: vec_data_103 = data_d1[255:248];
        7'd33: vec_data_103 = data_d1[263:256];
        7'd34: vec_data_103 = data_d1[271:264];
        7'd35: vec_data_103 = data_d1[279:272];
        7'd36: vec_data_103 = data_d1[287:280];
        7'd37: vec_data_103 = data_d1[295:288];
        7'd38: vec_data_103 = data_d1[303:296];
        7'd39: vec_data_103 = data_d1[311:304];
        7'd40: vec_data_103 = data_d1[319:312];
        7'd41: vec_data_103 = data_d1[327:320];
        7'd42: vec_data_103 = data_d1[335:328];
        7'd43: vec_data_103 = data_d1[343:336];
        7'd44: vec_data_103 = data_d1[351:344];
        7'd45: vec_data_103 = data_d1[359:352];
        7'd46: vec_data_103 = data_d1[367:360];
        7'd47: vec_data_103 = data_d1[375:368];
        7'd48: vec_data_103 = data_d1[383:376];
        7'd49: vec_data_103 = data_d1[391:384];
        7'd50: vec_data_103 = data_d1[399:392];
        7'd51: vec_data_103 = data_d1[407:400];
        7'd52: vec_data_103 = data_d1[415:408];
        7'd53: vec_data_103 = data_d1[423:416];
        7'd54: vec_data_103 = data_d1[431:424];
        7'd55: vec_data_103 = data_d1[439:432];
        7'd56: vec_data_103 = data_d1[447:440];
        7'd57: vec_data_103 = data_d1[455:448];
        7'd58: vec_data_103 = data_d1[463:456];
        7'd59: vec_data_103 = data_d1[471:464];
        7'd60: vec_data_103 = data_d1[479:472];
        7'd61: vec_data_103 = data_d1[487:480];
        7'd62: vec_data_103 = data_d1[495:488];
        7'd63: vec_data_103 = data_d1[503:496];
        7'd64: vec_data_103 = data_d1[511:504];
        7'd65: vec_data_103 = data_d1[519:512];
        7'd66: vec_data_103 = data_d1[527:520];
        7'd67: vec_data_103 = data_d1[535:528];
        7'd68: vec_data_103 = data_d1[543:536];
        7'd69: vec_data_103 = data_d1[551:544];
        7'd70: vec_data_103 = data_d1[559:552];
        7'd71: vec_data_103 = data_d1[567:560];
        7'd72: vec_data_103 = data_d1[575:568];
        7'd73: vec_data_103 = data_d1[583:576];
        7'd74: vec_data_103 = data_d1[591:584];
        7'd75: vec_data_103 = data_d1[599:592];
        7'd76: vec_data_103 = data_d1[607:600];
        7'd77: vec_data_103 = data_d1[615:608];
        7'd78: vec_data_103 = data_d1[623:616];
        7'd79: vec_data_103 = data_d1[631:624];
        7'd80: vec_data_103 = data_d1[639:632];
        7'd81: vec_data_103 = data_d1[647:640];
        7'd82: vec_data_103 = data_d1[655:648];
        7'd83: vec_data_103 = data_d1[663:656];
        7'd84: vec_data_103 = data_d1[671:664];
        7'd85: vec_data_103 = data_d1[679:672];
        7'd86: vec_data_103 = data_d1[687:680];
        7'd87: vec_data_103 = data_d1[695:688];
        7'd88: vec_data_103 = data_d1[703:696];
        7'd89: vec_data_103 = data_d1[711:704];
        7'd90: vec_data_103 = data_d1[719:712];
        7'd91: vec_data_103 = data_d1[727:720];
        7'd92: vec_data_103 = data_d1[735:728];
        7'd93: vec_data_103 = data_d1[743:736];
        7'd94: vec_data_103 = data_d1[751:744];
        7'd95: vec_data_103 = data_d1[759:752];
        7'd96: vec_data_103 = data_d1[767:760];
        7'd97: vec_data_103 = data_d1[775:768];
        7'd98: vec_data_103 = data_d1[783:776];
        7'd99: vec_data_103 = data_d1[791:784];
        7'd100: vec_data_103 = data_d1[799:792];
        7'd101: vec_data_103 = data_d1[807:800];
        7'd102: vec_data_103 = data_d1[815:808];
        7'd103: vec_data_103 = data_d1[823:816];
        7'd104: vec_data_103 = data_d1[831:824];
    endcase
end

always @(
  vec_sum_104_d1
  or data_d1
  ) begin
    vec_data_104 = 8'b0;
    case(vec_sum_104_d1)
        7'd1: vec_data_104 = data_d1[7:0];
        7'd2: vec_data_104 = data_d1[15:8];
        7'd3: vec_data_104 = data_d1[23:16];
        7'd4: vec_data_104 = data_d1[31:24];
        7'd5: vec_data_104 = data_d1[39:32];
        7'd6: vec_data_104 = data_d1[47:40];
        7'd7: vec_data_104 = data_d1[55:48];
        7'd8: vec_data_104 = data_d1[63:56];
        7'd9: vec_data_104 = data_d1[71:64];
        7'd10: vec_data_104 = data_d1[79:72];
        7'd11: vec_data_104 = data_d1[87:80];
        7'd12: vec_data_104 = data_d1[95:88];
        7'd13: vec_data_104 = data_d1[103:96];
        7'd14: vec_data_104 = data_d1[111:104];
        7'd15: vec_data_104 = data_d1[119:112];
        7'd16: vec_data_104 = data_d1[127:120];
        7'd17: vec_data_104 = data_d1[135:128];
        7'd18: vec_data_104 = data_d1[143:136];
        7'd19: vec_data_104 = data_d1[151:144];
        7'd20: vec_data_104 = data_d1[159:152];
        7'd21: vec_data_104 = data_d1[167:160];
        7'd22: vec_data_104 = data_d1[175:168];
        7'd23: vec_data_104 = data_d1[183:176];
        7'd24: vec_data_104 = data_d1[191:184];
        7'd25: vec_data_104 = data_d1[199:192];
        7'd26: vec_data_104 = data_d1[207:200];
        7'd27: vec_data_104 = data_d1[215:208];
        7'd28: vec_data_104 = data_d1[223:216];
        7'd29: vec_data_104 = data_d1[231:224];
        7'd30: vec_data_104 = data_d1[239:232];
        7'd31: vec_data_104 = data_d1[247:240];
        7'd32: vec_data_104 = data_d1[255:248];
        7'd33: vec_data_104 = data_d1[263:256];
        7'd34: vec_data_104 = data_d1[271:264];
        7'd35: vec_data_104 = data_d1[279:272];
        7'd36: vec_data_104 = data_d1[287:280];
        7'd37: vec_data_104 = data_d1[295:288];
        7'd38: vec_data_104 = data_d1[303:296];
        7'd39: vec_data_104 = data_d1[311:304];
        7'd40: vec_data_104 = data_d1[319:312];
        7'd41: vec_data_104 = data_d1[327:320];
        7'd42: vec_data_104 = data_d1[335:328];
        7'd43: vec_data_104 = data_d1[343:336];
        7'd44: vec_data_104 = data_d1[351:344];
        7'd45: vec_data_104 = data_d1[359:352];
        7'd46: vec_data_104 = data_d1[367:360];
        7'd47: vec_data_104 = data_d1[375:368];
        7'd48: vec_data_104 = data_d1[383:376];
        7'd49: vec_data_104 = data_d1[391:384];
        7'd50: vec_data_104 = data_d1[399:392];
        7'd51: vec_data_104 = data_d1[407:400];
        7'd52: vec_data_104 = data_d1[415:408];
        7'd53: vec_data_104 = data_d1[423:416];
        7'd54: vec_data_104 = data_d1[431:424];
        7'd55: vec_data_104 = data_d1[439:432];
        7'd56: vec_data_104 = data_d1[447:440];
        7'd57: vec_data_104 = data_d1[455:448];
        7'd58: vec_data_104 = data_d1[463:456];
        7'd59: vec_data_104 = data_d1[471:464];
        7'd60: vec_data_104 = data_d1[479:472];
        7'd61: vec_data_104 = data_d1[487:480];
        7'd62: vec_data_104 = data_d1[495:488];
        7'd63: vec_data_104 = data_d1[503:496];
        7'd64: vec_data_104 = data_d1[511:504];
        7'd65: vec_data_104 = data_d1[519:512];
        7'd66: vec_data_104 = data_d1[527:520];
        7'd67: vec_data_104 = data_d1[535:528];
        7'd68: vec_data_104 = data_d1[543:536];
        7'd69: vec_data_104 = data_d1[551:544];
        7'd70: vec_data_104 = data_d1[559:552];
        7'd71: vec_data_104 = data_d1[567:560];
        7'd72: vec_data_104 = data_d1[575:568];
        7'd73: vec_data_104 = data_d1[583:576];
        7'd74: vec_data_104 = data_d1[591:584];
        7'd75: vec_data_104 = data_d1[599:592];
        7'd76: vec_data_104 = data_d1[607:600];
        7'd77: vec_data_104 = data_d1[615:608];
        7'd78: vec_data_104 = data_d1[623:616];
        7'd79: vec_data_104 = data_d1[631:624];
        7'd80: vec_data_104 = data_d1[639:632];
        7'd81: vec_data_104 = data_d1[647:640];
        7'd82: vec_data_104 = data_d1[655:648];
        7'd83: vec_data_104 = data_d1[663:656];
        7'd84: vec_data_104 = data_d1[671:664];
        7'd85: vec_data_104 = data_d1[679:672];
        7'd86: vec_data_104 = data_d1[687:680];
        7'd87: vec_data_104 = data_d1[695:688];
        7'd88: vec_data_104 = data_d1[703:696];
        7'd89: vec_data_104 = data_d1[711:704];
        7'd90: vec_data_104 = data_d1[719:712];
        7'd91: vec_data_104 = data_d1[727:720];
        7'd92: vec_data_104 = data_d1[735:728];
        7'd93: vec_data_104 = data_d1[743:736];
        7'd94: vec_data_104 = data_d1[751:744];
        7'd95: vec_data_104 = data_d1[759:752];
        7'd96: vec_data_104 = data_d1[767:760];
        7'd97: vec_data_104 = data_d1[775:768];
        7'd98: vec_data_104 = data_d1[783:776];
        7'd99: vec_data_104 = data_d1[791:784];
        7'd100: vec_data_104 = data_d1[799:792];
        7'd101: vec_data_104 = data_d1[807:800];
        7'd102: vec_data_104 = data_d1[815:808];
        7'd103: vec_data_104 = data_d1[823:816];
        7'd104: vec_data_104 = data_d1[831:824];
        7'd105: vec_data_104 = data_d1[839:832];
    endcase
end

always @(
  vec_sum_105_d1
  or data_d1
  ) begin
    vec_data_105 = 8'b0;
    case(vec_sum_105_d1)
        7'd1: vec_data_105 = data_d1[7:0];
        7'd2: vec_data_105 = data_d1[15:8];
        7'd3: vec_data_105 = data_d1[23:16];
        7'd4: vec_data_105 = data_d1[31:24];
        7'd5: vec_data_105 = data_d1[39:32];
        7'd6: vec_data_105 = data_d1[47:40];
        7'd7: vec_data_105 = data_d1[55:48];
        7'd8: vec_data_105 = data_d1[63:56];
        7'd9: vec_data_105 = data_d1[71:64];
        7'd10: vec_data_105 = data_d1[79:72];
        7'd11: vec_data_105 = data_d1[87:80];
        7'd12: vec_data_105 = data_d1[95:88];
        7'd13: vec_data_105 = data_d1[103:96];
        7'd14: vec_data_105 = data_d1[111:104];
        7'd15: vec_data_105 = data_d1[119:112];
        7'd16: vec_data_105 = data_d1[127:120];
        7'd17: vec_data_105 = data_d1[135:128];
        7'd18: vec_data_105 = data_d1[143:136];
        7'd19: vec_data_105 = data_d1[151:144];
        7'd20: vec_data_105 = data_d1[159:152];
        7'd21: vec_data_105 = data_d1[167:160];
        7'd22: vec_data_105 = data_d1[175:168];
        7'd23: vec_data_105 = data_d1[183:176];
        7'd24: vec_data_105 = data_d1[191:184];
        7'd25: vec_data_105 = data_d1[199:192];
        7'd26: vec_data_105 = data_d1[207:200];
        7'd27: vec_data_105 = data_d1[215:208];
        7'd28: vec_data_105 = data_d1[223:216];
        7'd29: vec_data_105 = data_d1[231:224];
        7'd30: vec_data_105 = data_d1[239:232];
        7'd31: vec_data_105 = data_d1[247:240];
        7'd32: vec_data_105 = data_d1[255:248];
        7'd33: vec_data_105 = data_d1[263:256];
        7'd34: vec_data_105 = data_d1[271:264];
        7'd35: vec_data_105 = data_d1[279:272];
        7'd36: vec_data_105 = data_d1[287:280];
        7'd37: vec_data_105 = data_d1[295:288];
        7'd38: vec_data_105 = data_d1[303:296];
        7'd39: vec_data_105 = data_d1[311:304];
        7'd40: vec_data_105 = data_d1[319:312];
        7'd41: vec_data_105 = data_d1[327:320];
        7'd42: vec_data_105 = data_d1[335:328];
        7'd43: vec_data_105 = data_d1[343:336];
        7'd44: vec_data_105 = data_d1[351:344];
        7'd45: vec_data_105 = data_d1[359:352];
        7'd46: vec_data_105 = data_d1[367:360];
        7'd47: vec_data_105 = data_d1[375:368];
        7'd48: vec_data_105 = data_d1[383:376];
        7'd49: vec_data_105 = data_d1[391:384];
        7'd50: vec_data_105 = data_d1[399:392];
        7'd51: vec_data_105 = data_d1[407:400];
        7'd52: vec_data_105 = data_d1[415:408];
        7'd53: vec_data_105 = data_d1[423:416];
        7'd54: vec_data_105 = data_d1[431:424];
        7'd55: vec_data_105 = data_d1[439:432];
        7'd56: vec_data_105 = data_d1[447:440];
        7'd57: vec_data_105 = data_d1[455:448];
        7'd58: vec_data_105 = data_d1[463:456];
        7'd59: vec_data_105 = data_d1[471:464];
        7'd60: vec_data_105 = data_d1[479:472];
        7'd61: vec_data_105 = data_d1[487:480];
        7'd62: vec_data_105 = data_d1[495:488];
        7'd63: vec_data_105 = data_d1[503:496];
        7'd64: vec_data_105 = data_d1[511:504];
        7'd65: vec_data_105 = data_d1[519:512];
        7'd66: vec_data_105 = data_d1[527:520];
        7'd67: vec_data_105 = data_d1[535:528];
        7'd68: vec_data_105 = data_d1[543:536];
        7'd69: vec_data_105 = data_d1[551:544];
        7'd70: vec_data_105 = data_d1[559:552];
        7'd71: vec_data_105 = data_d1[567:560];
        7'd72: vec_data_105 = data_d1[575:568];
        7'd73: vec_data_105 = data_d1[583:576];
        7'd74: vec_data_105 = data_d1[591:584];
        7'd75: vec_data_105 = data_d1[599:592];
        7'd76: vec_data_105 = data_d1[607:600];
        7'd77: vec_data_105 = data_d1[615:608];
        7'd78: vec_data_105 = data_d1[623:616];
        7'd79: vec_data_105 = data_d1[631:624];
        7'd80: vec_data_105 = data_d1[639:632];
        7'd81: vec_data_105 = data_d1[647:640];
        7'd82: vec_data_105 = data_d1[655:648];
        7'd83: vec_data_105 = data_d1[663:656];
        7'd84: vec_data_105 = data_d1[671:664];
        7'd85: vec_data_105 = data_d1[679:672];
        7'd86: vec_data_105 = data_d1[687:680];
        7'd87: vec_data_105 = data_d1[695:688];
        7'd88: vec_data_105 = data_d1[703:696];
        7'd89: vec_data_105 = data_d1[711:704];
        7'd90: vec_data_105 = data_d1[719:712];
        7'd91: vec_data_105 = data_d1[727:720];
        7'd92: vec_data_105 = data_d1[735:728];
        7'd93: vec_data_105 = data_d1[743:736];
        7'd94: vec_data_105 = data_d1[751:744];
        7'd95: vec_data_105 = data_d1[759:752];
        7'd96: vec_data_105 = data_d1[767:760];
        7'd97: vec_data_105 = data_d1[775:768];
        7'd98: vec_data_105 = data_d1[783:776];
        7'd99: vec_data_105 = data_d1[791:784];
        7'd100: vec_data_105 = data_d1[799:792];
        7'd101: vec_data_105 = data_d1[807:800];
        7'd102: vec_data_105 = data_d1[815:808];
        7'd103: vec_data_105 = data_d1[823:816];
        7'd104: vec_data_105 = data_d1[831:824];
        7'd105: vec_data_105 = data_d1[839:832];
        7'd106: vec_data_105 = data_d1[847:840];
    endcase
end

always @(
  vec_sum_106_d1
  or data_d1
  ) begin
    vec_data_106 = 8'b0;
    case(vec_sum_106_d1)
        7'd1: vec_data_106 = data_d1[7:0];
        7'd2: vec_data_106 = data_d1[15:8];
        7'd3: vec_data_106 = data_d1[23:16];
        7'd4: vec_data_106 = data_d1[31:24];
        7'd5: vec_data_106 = data_d1[39:32];
        7'd6: vec_data_106 = data_d1[47:40];
        7'd7: vec_data_106 = data_d1[55:48];
        7'd8: vec_data_106 = data_d1[63:56];
        7'd9: vec_data_106 = data_d1[71:64];
        7'd10: vec_data_106 = data_d1[79:72];
        7'd11: vec_data_106 = data_d1[87:80];
        7'd12: vec_data_106 = data_d1[95:88];
        7'd13: vec_data_106 = data_d1[103:96];
        7'd14: vec_data_106 = data_d1[111:104];
        7'd15: vec_data_106 = data_d1[119:112];
        7'd16: vec_data_106 = data_d1[127:120];
        7'd17: vec_data_106 = data_d1[135:128];
        7'd18: vec_data_106 = data_d1[143:136];
        7'd19: vec_data_106 = data_d1[151:144];
        7'd20: vec_data_106 = data_d1[159:152];
        7'd21: vec_data_106 = data_d1[167:160];
        7'd22: vec_data_106 = data_d1[175:168];
        7'd23: vec_data_106 = data_d1[183:176];
        7'd24: vec_data_106 = data_d1[191:184];
        7'd25: vec_data_106 = data_d1[199:192];
        7'd26: vec_data_106 = data_d1[207:200];
        7'd27: vec_data_106 = data_d1[215:208];
        7'd28: vec_data_106 = data_d1[223:216];
        7'd29: vec_data_106 = data_d1[231:224];
        7'd30: vec_data_106 = data_d1[239:232];
        7'd31: vec_data_106 = data_d1[247:240];
        7'd32: vec_data_106 = data_d1[255:248];
        7'd33: vec_data_106 = data_d1[263:256];
        7'd34: vec_data_106 = data_d1[271:264];
        7'd35: vec_data_106 = data_d1[279:272];
        7'd36: vec_data_106 = data_d1[287:280];
        7'd37: vec_data_106 = data_d1[295:288];
        7'd38: vec_data_106 = data_d1[303:296];
        7'd39: vec_data_106 = data_d1[311:304];
        7'd40: vec_data_106 = data_d1[319:312];
        7'd41: vec_data_106 = data_d1[327:320];
        7'd42: vec_data_106 = data_d1[335:328];
        7'd43: vec_data_106 = data_d1[343:336];
        7'd44: vec_data_106 = data_d1[351:344];
        7'd45: vec_data_106 = data_d1[359:352];
        7'd46: vec_data_106 = data_d1[367:360];
        7'd47: vec_data_106 = data_d1[375:368];
        7'd48: vec_data_106 = data_d1[383:376];
        7'd49: vec_data_106 = data_d1[391:384];
        7'd50: vec_data_106 = data_d1[399:392];
        7'd51: vec_data_106 = data_d1[407:400];
        7'd52: vec_data_106 = data_d1[415:408];
        7'd53: vec_data_106 = data_d1[423:416];
        7'd54: vec_data_106 = data_d1[431:424];
        7'd55: vec_data_106 = data_d1[439:432];
        7'd56: vec_data_106 = data_d1[447:440];
        7'd57: vec_data_106 = data_d1[455:448];
        7'd58: vec_data_106 = data_d1[463:456];
        7'd59: vec_data_106 = data_d1[471:464];
        7'd60: vec_data_106 = data_d1[479:472];
        7'd61: vec_data_106 = data_d1[487:480];
        7'd62: vec_data_106 = data_d1[495:488];
        7'd63: vec_data_106 = data_d1[503:496];
        7'd64: vec_data_106 = data_d1[511:504];
        7'd65: vec_data_106 = data_d1[519:512];
        7'd66: vec_data_106 = data_d1[527:520];
        7'd67: vec_data_106 = data_d1[535:528];
        7'd68: vec_data_106 = data_d1[543:536];
        7'd69: vec_data_106 = data_d1[551:544];
        7'd70: vec_data_106 = data_d1[559:552];
        7'd71: vec_data_106 = data_d1[567:560];
        7'd72: vec_data_106 = data_d1[575:568];
        7'd73: vec_data_106 = data_d1[583:576];
        7'd74: vec_data_106 = data_d1[591:584];
        7'd75: vec_data_106 = data_d1[599:592];
        7'd76: vec_data_106 = data_d1[607:600];
        7'd77: vec_data_106 = data_d1[615:608];
        7'd78: vec_data_106 = data_d1[623:616];
        7'd79: vec_data_106 = data_d1[631:624];
        7'd80: vec_data_106 = data_d1[639:632];
        7'd81: vec_data_106 = data_d1[647:640];
        7'd82: vec_data_106 = data_d1[655:648];
        7'd83: vec_data_106 = data_d1[663:656];
        7'd84: vec_data_106 = data_d1[671:664];
        7'd85: vec_data_106 = data_d1[679:672];
        7'd86: vec_data_106 = data_d1[687:680];
        7'd87: vec_data_106 = data_d1[695:688];
        7'd88: vec_data_106 = data_d1[703:696];
        7'd89: vec_data_106 = data_d1[711:704];
        7'd90: vec_data_106 = data_d1[719:712];
        7'd91: vec_data_106 = data_d1[727:720];
        7'd92: vec_data_106 = data_d1[735:728];
        7'd93: vec_data_106 = data_d1[743:736];
        7'd94: vec_data_106 = data_d1[751:744];
        7'd95: vec_data_106 = data_d1[759:752];
        7'd96: vec_data_106 = data_d1[767:760];
        7'd97: vec_data_106 = data_d1[775:768];
        7'd98: vec_data_106 = data_d1[783:776];
        7'd99: vec_data_106 = data_d1[791:784];
        7'd100: vec_data_106 = data_d1[799:792];
        7'd101: vec_data_106 = data_d1[807:800];
        7'd102: vec_data_106 = data_d1[815:808];
        7'd103: vec_data_106 = data_d1[823:816];
        7'd104: vec_data_106 = data_d1[831:824];
        7'd105: vec_data_106 = data_d1[839:832];
        7'd106: vec_data_106 = data_d1[847:840];
        7'd107: vec_data_106 = data_d1[855:848];
    endcase
end

always @(
  vec_sum_107_d1
  or data_d1
  ) begin
    vec_data_107 = 8'b0;
    case(vec_sum_107_d1)
        7'd1: vec_data_107 = data_d1[7:0];
        7'd2: vec_data_107 = data_d1[15:8];
        7'd3: vec_data_107 = data_d1[23:16];
        7'd4: vec_data_107 = data_d1[31:24];
        7'd5: vec_data_107 = data_d1[39:32];
        7'd6: vec_data_107 = data_d1[47:40];
        7'd7: vec_data_107 = data_d1[55:48];
        7'd8: vec_data_107 = data_d1[63:56];
        7'd9: vec_data_107 = data_d1[71:64];
        7'd10: vec_data_107 = data_d1[79:72];
        7'd11: vec_data_107 = data_d1[87:80];
        7'd12: vec_data_107 = data_d1[95:88];
        7'd13: vec_data_107 = data_d1[103:96];
        7'd14: vec_data_107 = data_d1[111:104];
        7'd15: vec_data_107 = data_d1[119:112];
        7'd16: vec_data_107 = data_d1[127:120];
        7'd17: vec_data_107 = data_d1[135:128];
        7'd18: vec_data_107 = data_d1[143:136];
        7'd19: vec_data_107 = data_d1[151:144];
        7'd20: vec_data_107 = data_d1[159:152];
        7'd21: vec_data_107 = data_d1[167:160];
        7'd22: vec_data_107 = data_d1[175:168];
        7'd23: vec_data_107 = data_d1[183:176];
        7'd24: vec_data_107 = data_d1[191:184];
        7'd25: vec_data_107 = data_d1[199:192];
        7'd26: vec_data_107 = data_d1[207:200];
        7'd27: vec_data_107 = data_d1[215:208];
        7'd28: vec_data_107 = data_d1[223:216];
        7'd29: vec_data_107 = data_d1[231:224];
        7'd30: vec_data_107 = data_d1[239:232];
        7'd31: vec_data_107 = data_d1[247:240];
        7'd32: vec_data_107 = data_d1[255:248];
        7'd33: vec_data_107 = data_d1[263:256];
        7'd34: vec_data_107 = data_d1[271:264];
        7'd35: vec_data_107 = data_d1[279:272];
        7'd36: vec_data_107 = data_d1[287:280];
        7'd37: vec_data_107 = data_d1[295:288];
        7'd38: vec_data_107 = data_d1[303:296];
        7'd39: vec_data_107 = data_d1[311:304];
        7'd40: vec_data_107 = data_d1[319:312];
        7'd41: vec_data_107 = data_d1[327:320];
        7'd42: vec_data_107 = data_d1[335:328];
        7'd43: vec_data_107 = data_d1[343:336];
        7'd44: vec_data_107 = data_d1[351:344];
        7'd45: vec_data_107 = data_d1[359:352];
        7'd46: vec_data_107 = data_d1[367:360];
        7'd47: vec_data_107 = data_d1[375:368];
        7'd48: vec_data_107 = data_d1[383:376];
        7'd49: vec_data_107 = data_d1[391:384];
        7'd50: vec_data_107 = data_d1[399:392];
        7'd51: vec_data_107 = data_d1[407:400];
        7'd52: vec_data_107 = data_d1[415:408];
        7'd53: vec_data_107 = data_d1[423:416];
        7'd54: vec_data_107 = data_d1[431:424];
        7'd55: vec_data_107 = data_d1[439:432];
        7'd56: vec_data_107 = data_d1[447:440];
        7'd57: vec_data_107 = data_d1[455:448];
        7'd58: vec_data_107 = data_d1[463:456];
        7'd59: vec_data_107 = data_d1[471:464];
        7'd60: vec_data_107 = data_d1[479:472];
        7'd61: vec_data_107 = data_d1[487:480];
        7'd62: vec_data_107 = data_d1[495:488];
        7'd63: vec_data_107 = data_d1[503:496];
        7'd64: vec_data_107 = data_d1[511:504];
        7'd65: vec_data_107 = data_d1[519:512];
        7'd66: vec_data_107 = data_d1[527:520];
        7'd67: vec_data_107 = data_d1[535:528];
        7'd68: vec_data_107 = data_d1[543:536];
        7'd69: vec_data_107 = data_d1[551:544];
        7'd70: vec_data_107 = data_d1[559:552];
        7'd71: vec_data_107 = data_d1[567:560];
        7'd72: vec_data_107 = data_d1[575:568];
        7'd73: vec_data_107 = data_d1[583:576];
        7'd74: vec_data_107 = data_d1[591:584];
        7'd75: vec_data_107 = data_d1[599:592];
        7'd76: vec_data_107 = data_d1[607:600];
        7'd77: vec_data_107 = data_d1[615:608];
        7'd78: vec_data_107 = data_d1[623:616];
        7'd79: vec_data_107 = data_d1[631:624];
        7'd80: vec_data_107 = data_d1[639:632];
        7'd81: vec_data_107 = data_d1[647:640];
        7'd82: vec_data_107 = data_d1[655:648];
        7'd83: vec_data_107 = data_d1[663:656];
        7'd84: vec_data_107 = data_d1[671:664];
        7'd85: vec_data_107 = data_d1[679:672];
        7'd86: vec_data_107 = data_d1[687:680];
        7'd87: vec_data_107 = data_d1[695:688];
        7'd88: vec_data_107 = data_d1[703:696];
        7'd89: vec_data_107 = data_d1[711:704];
        7'd90: vec_data_107 = data_d1[719:712];
        7'd91: vec_data_107 = data_d1[727:720];
        7'd92: vec_data_107 = data_d1[735:728];
        7'd93: vec_data_107 = data_d1[743:736];
        7'd94: vec_data_107 = data_d1[751:744];
        7'd95: vec_data_107 = data_d1[759:752];
        7'd96: vec_data_107 = data_d1[767:760];
        7'd97: vec_data_107 = data_d1[775:768];
        7'd98: vec_data_107 = data_d1[783:776];
        7'd99: vec_data_107 = data_d1[791:784];
        7'd100: vec_data_107 = data_d1[799:792];
        7'd101: vec_data_107 = data_d1[807:800];
        7'd102: vec_data_107 = data_d1[815:808];
        7'd103: vec_data_107 = data_d1[823:816];
        7'd104: vec_data_107 = data_d1[831:824];
        7'd105: vec_data_107 = data_d1[839:832];
        7'd106: vec_data_107 = data_d1[847:840];
        7'd107: vec_data_107 = data_d1[855:848];
        7'd108: vec_data_107 = data_d1[863:856];
    endcase
end

always @(
  vec_sum_108_d1
  or data_d1
  ) begin
    vec_data_108 = 8'b0;
    case(vec_sum_108_d1)
        7'd1: vec_data_108 = data_d1[7:0];
        7'd2: vec_data_108 = data_d1[15:8];
        7'd3: vec_data_108 = data_d1[23:16];
        7'd4: vec_data_108 = data_d1[31:24];
        7'd5: vec_data_108 = data_d1[39:32];
        7'd6: vec_data_108 = data_d1[47:40];
        7'd7: vec_data_108 = data_d1[55:48];
        7'd8: vec_data_108 = data_d1[63:56];
        7'd9: vec_data_108 = data_d1[71:64];
        7'd10: vec_data_108 = data_d1[79:72];
        7'd11: vec_data_108 = data_d1[87:80];
        7'd12: vec_data_108 = data_d1[95:88];
        7'd13: vec_data_108 = data_d1[103:96];
        7'd14: vec_data_108 = data_d1[111:104];
        7'd15: vec_data_108 = data_d1[119:112];
        7'd16: vec_data_108 = data_d1[127:120];
        7'd17: vec_data_108 = data_d1[135:128];
        7'd18: vec_data_108 = data_d1[143:136];
        7'd19: vec_data_108 = data_d1[151:144];
        7'd20: vec_data_108 = data_d1[159:152];
        7'd21: vec_data_108 = data_d1[167:160];
        7'd22: vec_data_108 = data_d1[175:168];
        7'd23: vec_data_108 = data_d1[183:176];
        7'd24: vec_data_108 = data_d1[191:184];
        7'd25: vec_data_108 = data_d1[199:192];
        7'd26: vec_data_108 = data_d1[207:200];
        7'd27: vec_data_108 = data_d1[215:208];
        7'd28: vec_data_108 = data_d1[223:216];
        7'd29: vec_data_108 = data_d1[231:224];
        7'd30: vec_data_108 = data_d1[239:232];
        7'd31: vec_data_108 = data_d1[247:240];
        7'd32: vec_data_108 = data_d1[255:248];
        7'd33: vec_data_108 = data_d1[263:256];
        7'd34: vec_data_108 = data_d1[271:264];
        7'd35: vec_data_108 = data_d1[279:272];
        7'd36: vec_data_108 = data_d1[287:280];
        7'd37: vec_data_108 = data_d1[295:288];
        7'd38: vec_data_108 = data_d1[303:296];
        7'd39: vec_data_108 = data_d1[311:304];
        7'd40: vec_data_108 = data_d1[319:312];
        7'd41: vec_data_108 = data_d1[327:320];
        7'd42: vec_data_108 = data_d1[335:328];
        7'd43: vec_data_108 = data_d1[343:336];
        7'd44: vec_data_108 = data_d1[351:344];
        7'd45: vec_data_108 = data_d1[359:352];
        7'd46: vec_data_108 = data_d1[367:360];
        7'd47: vec_data_108 = data_d1[375:368];
        7'd48: vec_data_108 = data_d1[383:376];
        7'd49: vec_data_108 = data_d1[391:384];
        7'd50: vec_data_108 = data_d1[399:392];
        7'd51: vec_data_108 = data_d1[407:400];
        7'd52: vec_data_108 = data_d1[415:408];
        7'd53: vec_data_108 = data_d1[423:416];
        7'd54: vec_data_108 = data_d1[431:424];
        7'd55: vec_data_108 = data_d1[439:432];
        7'd56: vec_data_108 = data_d1[447:440];
        7'd57: vec_data_108 = data_d1[455:448];
        7'd58: vec_data_108 = data_d1[463:456];
        7'd59: vec_data_108 = data_d1[471:464];
        7'd60: vec_data_108 = data_d1[479:472];
        7'd61: vec_data_108 = data_d1[487:480];
        7'd62: vec_data_108 = data_d1[495:488];
        7'd63: vec_data_108 = data_d1[503:496];
        7'd64: vec_data_108 = data_d1[511:504];
        7'd65: vec_data_108 = data_d1[519:512];
        7'd66: vec_data_108 = data_d1[527:520];
        7'd67: vec_data_108 = data_d1[535:528];
        7'd68: vec_data_108 = data_d1[543:536];
        7'd69: vec_data_108 = data_d1[551:544];
        7'd70: vec_data_108 = data_d1[559:552];
        7'd71: vec_data_108 = data_d1[567:560];
        7'd72: vec_data_108 = data_d1[575:568];
        7'd73: vec_data_108 = data_d1[583:576];
        7'd74: vec_data_108 = data_d1[591:584];
        7'd75: vec_data_108 = data_d1[599:592];
        7'd76: vec_data_108 = data_d1[607:600];
        7'd77: vec_data_108 = data_d1[615:608];
        7'd78: vec_data_108 = data_d1[623:616];
        7'd79: vec_data_108 = data_d1[631:624];
        7'd80: vec_data_108 = data_d1[639:632];
        7'd81: vec_data_108 = data_d1[647:640];
        7'd82: vec_data_108 = data_d1[655:648];
        7'd83: vec_data_108 = data_d1[663:656];
        7'd84: vec_data_108 = data_d1[671:664];
        7'd85: vec_data_108 = data_d1[679:672];
        7'd86: vec_data_108 = data_d1[687:680];
        7'd87: vec_data_108 = data_d1[695:688];
        7'd88: vec_data_108 = data_d1[703:696];
        7'd89: vec_data_108 = data_d1[711:704];
        7'd90: vec_data_108 = data_d1[719:712];
        7'd91: vec_data_108 = data_d1[727:720];
        7'd92: vec_data_108 = data_d1[735:728];
        7'd93: vec_data_108 = data_d1[743:736];
        7'd94: vec_data_108 = data_d1[751:744];
        7'd95: vec_data_108 = data_d1[759:752];
        7'd96: vec_data_108 = data_d1[767:760];
        7'd97: vec_data_108 = data_d1[775:768];
        7'd98: vec_data_108 = data_d1[783:776];
        7'd99: vec_data_108 = data_d1[791:784];
        7'd100: vec_data_108 = data_d1[799:792];
        7'd101: vec_data_108 = data_d1[807:800];
        7'd102: vec_data_108 = data_d1[815:808];
        7'd103: vec_data_108 = data_d1[823:816];
        7'd104: vec_data_108 = data_d1[831:824];
        7'd105: vec_data_108 = data_d1[839:832];
        7'd106: vec_data_108 = data_d1[847:840];
        7'd107: vec_data_108 = data_d1[855:848];
        7'd108: vec_data_108 = data_d1[863:856];
        7'd109: vec_data_108 = data_d1[871:864];
    endcase
end

always @(
  vec_sum_109_d1
  or data_d1
  ) begin
    vec_data_109 = 8'b0;
    case(vec_sum_109_d1)
        7'd1: vec_data_109 = data_d1[7:0];
        7'd2: vec_data_109 = data_d1[15:8];
        7'd3: vec_data_109 = data_d1[23:16];
        7'd4: vec_data_109 = data_d1[31:24];
        7'd5: vec_data_109 = data_d1[39:32];
        7'd6: vec_data_109 = data_d1[47:40];
        7'd7: vec_data_109 = data_d1[55:48];
        7'd8: vec_data_109 = data_d1[63:56];
        7'd9: vec_data_109 = data_d1[71:64];
        7'd10: vec_data_109 = data_d1[79:72];
        7'd11: vec_data_109 = data_d1[87:80];
        7'd12: vec_data_109 = data_d1[95:88];
        7'd13: vec_data_109 = data_d1[103:96];
        7'd14: vec_data_109 = data_d1[111:104];
        7'd15: vec_data_109 = data_d1[119:112];
        7'd16: vec_data_109 = data_d1[127:120];
        7'd17: vec_data_109 = data_d1[135:128];
        7'd18: vec_data_109 = data_d1[143:136];
        7'd19: vec_data_109 = data_d1[151:144];
        7'd20: vec_data_109 = data_d1[159:152];
        7'd21: vec_data_109 = data_d1[167:160];
        7'd22: vec_data_109 = data_d1[175:168];
        7'd23: vec_data_109 = data_d1[183:176];
        7'd24: vec_data_109 = data_d1[191:184];
        7'd25: vec_data_109 = data_d1[199:192];
        7'd26: vec_data_109 = data_d1[207:200];
        7'd27: vec_data_109 = data_d1[215:208];
        7'd28: vec_data_109 = data_d1[223:216];
        7'd29: vec_data_109 = data_d1[231:224];
        7'd30: vec_data_109 = data_d1[239:232];
        7'd31: vec_data_109 = data_d1[247:240];
        7'd32: vec_data_109 = data_d1[255:248];
        7'd33: vec_data_109 = data_d1[263:256];
        7'd34: vec_data_109 = data_d1[271:264];
        7'd35: vec_data_109 = data_d1[279:272];
        7'd36: vec_data_109 = data_d1[287:280];
        7'd37: vec_data_109 = data_d1[295:288];
        7'd38: vec_data_109 = data_d1[303:296];
        7'd39: vec_data_109 = data_d1[311:304];
        7'd40: vec_data_109 = data_d1[319:312];
        7'd41: vec_data_109 = data_d1[327:320];
        7'd42: vec_data_109 = data_d1[335:328];
        7'd43: vec_data_109 = data_d1[343:336];
        7'd44: vec_data_109 = data_d1[351:344];
        7'd45: vec_data_109 = data_d1[359:352];
        7'd46: vec_data_109 = data_d1[367:360];
        7'd47: vec_data_109 = data_d1[375:368];
        7'd48: vec_data_109 = data_d1[383:376];
        7'd49: vec_data_109 = data_d1[391:384];
        7'd50: vec_data_109 = data_d1[399:392];
        7'd51: vec_data_109 = data_d1[407:400];
        7'd52: vec_data_109 = data_d1[415:408];
        7'd53: vec_data_109 = data_d1[423:416];
        7'd54: vec_data_109 = data_d1[431:424];
        7'd55: vec_data_109 = data_d1[439:432];
        7'd56: vec_data_109 = data_d1[447:440];
        7'd57: vec_data_109 = data_d1[455:448];
        7'd58: vec_data_109 = data_d1[463:456];
        7'd59: vec_data_109 = data_d1[471:464];
        7'd60: vec_data_109 = data_d1[479:472];
        7'd61: vec_data_109 = data_d1[487:480];
        7'd62: vec_data_109 = data_d1[495:488];
        7'd63: vec_data_109 = data_d1[503:496];
        7'd64: vec_data_109 = data_d1[511:504];
        7'd65: vec_data_109 = data_d1[519:512];
        7'd66: vec_data_109 = data_d1[527:520];
        7'd67: vec_data_109 = data_d1[535:528];
        7'd68: vec_data_109 = data_d1[543:536];
        7'd69: vec_data_109 = data_d1[551:544];
        7'd70: vec_data_109 = data_d1[559:552];
        7'd71: vec_data_109 = data_d1[567:560];
        7'd72: vec_data_109 = data_d1[575:568];
        7'd73: vec_data_109 = data_d1[583:576];
        7'd74: vec_data_109 = data_d1[591:584];
        7'd75: vec_data_109 = data_d1[599:592];
        7'd76: vec_data_109 = data_d1[607:600];
        7'd77: vec_data_109 = data_d1[615:608];
        7'd78: vec_data_109 = data_d1[623:616];
        7'd79: vec_data_109 = data_d1[631:624];
        7'd80: vec_data_109 = data_d1[639:632];
        7'd81: vec_data_109 = data_d1[647:640];
        7'd82: vec_data_109 = data_d1[655:648];
        7'd83: vec_data_109 = data_d1[663:656];
        7'd84: vec_data_109 = data_d1[671:664];
        7'd85: vec_data_109 = data_d1[679:672];
        7'd86: vec_data_109 = data_d1[687:680];
        7'd87: vec_data_109 = data_d1[695:688];
        7'd88: vec_data_109 = data_d1[703:696];
        7'd89: vec_data_109 = data_d1[711:704];
        7'd90: vec_data_109 = data_d1[719:712];
        7'd91: vec_data_109 = data_d1[727:720];
        7'd92: vec_data_109 = data_d1[735:728];
        7'd93: vec_data_109 = data_d1[743:736];
        7'd94: vec_data_109 = data_d1[751:744];
        7'd95: vec_data_109 = data_d1[759:752];
        7'd96: vec_data_109 = data_d1[767:760];
        7'd97: vec_data_109 = data_d1[775:768];
        7'd98: vec_data_109 = data_d1[783:776];
        7'd99: vec_data_109 = data_d1[791:784];
        7'd100: vec_data_109 = data_d1[799:792];
        7'd101: vec_data_109 = data_d1[807:800];
        7'd102: vec_data_109 = data_d1[815:808];
        7'd103: vec_data_109 = data_d1[823:816];
        7'd104: vec_data_109 = data_d1[831:824];
        7'd105: vec_data_109 = data_d1[839:832];
        7'd106: vec_data_109 = data_d1[847:840];
        7'd107: vec_data_109 = data_d1[855:848];
        7'd108: vec_data_109 = data_d1[863:856];
        7'd109: vec_data_109 = data_d1[871:864];
        7'd110: vec_data_109 = data_d1[879:872];
    endcase
end

always @(
  vec_sum_110_d1
  or data_d1
  ) begin
    vec_data_110 = 8'b0;
    case(vec_sum_110_d1)
        7'd1: vec_data_110 = data_d1[7:0];
        7'd2: vec_data_110 = data_d1[15:8];
        7'd3: vec_data_110 = data_d1[23:16];
        7'd4: vec_data_110 = data_d1[31:24];
        7'd5: vec_data_110 = data_d1[39:32];
        7'd6: vec_data_110 = data_d1[47:40];
        7'd7: vec_data_110 = data_d1[55:48];
        7'd8: vec_data_110 = data_d1[63:56];
        7'd9: vec_data_110 = data_d1[71:64];
        7'd10: vec_data_110 = data_d1[79:72];
        7'd11: vec_data_110 = data_d1[87:80];
        7'd12: vec_data_110 = data_d1[95:88];
        7'd13: vec_data_110 = data_d1[103:96];
        7'd14: vec_data_110 = data_d1[111:104];
        7'd15: vec_data_110 = data_d1[119:112];
        7'd16: vec_data_110 = data_d1[127:120];
        7'd17: vec_data_110 = data_d1[135:128];
        7'd18: vec_data_110 = data_d1[143:136];
        7'd19: vec_data_110 = data_d1[151:144];
        7'd20: vec_data_110 = data_d1[159:152];
        7'd21: vec_data_110 = data_d1[167:160];
        7'd22: vec_data_110 = data_d1[175:168];
        7'd23: vec_data_110 = data_d1[183:176];
        7'd24: vec_data_110 = data_d1[191:184];
        7'd25: vec_data_110 = data_d1[199:192];
        7'd26: vec_data_110 = data_d1[207:200];
        7'd27: vec_data_110 = data_d1[215:208];
        7'd28: vec_data_110 = data_d1[223:216];
        7'd29: vec_data_110 = data_d1[231:224];
        7'd30: vec_data_110 = data_d1[239:232];
        7'd31: vec_data_110 = data_d1[247:240];
        7'd32: vec_data_110 = data_d1[255:248];
        7'd33: vec_data_110 = data_d1[263:256];
        7'd34: vec_data_110 = data_d1[271:264];
        7'd35: vec_data_110 = data_d1[279:272];
        7'd36: vec_data_110 = data_d1[287:280];
        7'd37: vec_data_110 = data_d1[295:288];
        7'd38: vec_data_110 = data_d1[303:296];
        7'd39: vec_data_110 = data_d1[311:304];
        7'd40: vec_data_110 = data_d1[319:312];
        7'd41: vec_data_110 = data_d1[327:320];
        7'd42: vec_data_110 = data_d1[335:328];
        7'd43: vec_data_110 = data_d1[343:336];
        7'd44: vec_data_110 = data_d1[351:344];
        7'd45: vec_data_110 = data_d1[359:352];
        7'd46: vec_data_110 = data_d1[367:360];
        7'd47: vec_data_110 = data_d1[375:368];
        7'd48: vec_data_110 = data_d1[383:376];
        7'd49: vec_data_110 = data_d1[391:384];
        7'd50: vec_data_110 = data_d1[399:392];
        7'd51: vec_data_110 = data_d1[407:400];
        7'd52: vec_data_110 = data_d1[415:408];
        7'd53: vec_data_110 = data_d1[423:416];
        7'd54: vec_data_110 = data_d1[431:424];
        7'd55: vec_data_110 = data_d1[439:432];
        7'd56: vec_data_110 = data_d1[447:440];
        7'd57: vec_data_110 = data_d1[455:448];
        7'd58: vec_data_110 = data_d1[463:456];
        7'd59: vec_data_110 = data_d1[471:464];
        7'd60: vec_data_110 = data_d1[479:472];
        7'd61: vec_data_110 = data_d1[487:480];
        7'd62: vec_data_110 = data_d1[495:488];
        7'd63: vec_data_110 = data_d1[503:496];
        7'd64: vec_data_110 = data_d1[511:504];
        7'd65: vec_data_110 = data_d1[519:512];
        7'd66: vec_data_110 = data_d1[527:520];
        7'd67: vec_data_110 = data_d1[535:528];
        7'd68: vec_data_110 = data_d1[543:536];
        7'd69: vec_data_110 = data_d1[551:544];
        7'd70: vec_data_110 = data_d1[559:552];
        7'd71: vec_data_110 = data_d1[567:560];
        7'd72: vec_data_110 = data_d1[575:568];
        7'd73: vec_data_110 = data_d1[583:576];
        7'd74: vec_data_110 = data_d1[591:584];
        7'd75: vec_data_110 = data_d1[599:592];
        7'd76: vec_data_110 = data_d1[607:600];
        7'd77: vec_data_110 = data_d1[615:608];
        7'd78: vec_data_110 = data_d1[623:616];
        7'd79: vec_data_110 = data_d1[631:624];
        7'd80: vec_data_110 = data_d1[639:632];
        7'd81: vec_data_110 = data_d1[647:640];
        7'd82: vec_data_110 = data_d1[655:648];
        7'd83: vec_data_110 = data_d1[663:656];
        7'd84: vec_data_110 = data_d1[671:664];
        7'd85: vec_data_110 = data_d1[679:672];
        7'd86: vec_data_110 = data_d1[687:680];
        7'd87: vec_data_110 = data_d1[695:688];
        7'd88: vec_data_110 = data_d1[703:696];
        7'd89: vec_data_110 = data_d1[711:704];
        7'd90: vec_data_110 = data_d1[719:712];
        7'd91: vec_data_110 = data_d1[727:720];
        7'd92: vec_data_110 = data_d1[735:728];
        7'd93: vec_data_110 = data_d1[743:736];
        7'd94: vec_data_110 = data_d1[751:744];
        7'd95: vec_data_110 = data_d1[759:752];
        7'd96: vec_data_110 = data_d1[767:760];
        7'd97: vec_data_110 = data_d1[775:768];
        7'd98: vec_data_110 = data_d1[783:776];
        7'd99: vec_data_110 = data_d1[791:784];
        7'd100: vec_data_110 = data_d1[799:792];
        7'd101: vec_data_110 = data_d1[807:800];
        7'd102: vec_data_110 = data_d1[815:808];
        7'd103: vec_data_110 = data_d1[823:816];
        7'd104: vec_data_110 = data_d1[831:824];
        7'd105: vec_data_110 = data_d1[839:832];
        7'd106: vec_data_110 = data_d1[847:840];
        7'd107: vec_data_110 = data_d1[855:848];
        7'd108: vec_data_110 = data_d1[863:856];
        7'd109: vec_data_110 = data_d1[871:864];
        7'd110: vec_data_110 = data_d1[879:872];
        7'd111: vec_data_110 = data_d1[887:880];
    endcase
end

always @(
  vec_sum_111_d1
  or data_d1
  ) begin
    vec_data_111 = 8'b0;
    case(vec_sum_111_d1)
        7'd1: vec_data_111 = data_d1[7:0];
        7'd2: vec_data_111 = data_d1[15:8];
        7'd3: vec_data_111 = data_d1[23:16];
        7'd4: vec_data_111 = data_d1[31:24];
        7'd5: vec_data_111 = data_d1[39:32];
        7'd6: vec_data_111 = data_d1[47:40];
        7'd7: vec_data_111 = data_d1[55:48];
        7'd8: vec_data_111 = data_d1[63:56];
        7'd9: vec_data_111 = data_d1[71:64];
        7'd10: vec_data_111 = data_d1[79:72];
        7'd11: vec_data_111 = data_d1[87:80];
        7'd12: vec_data_111 = data_d1[95:88];
        7'd13: vec_data_111 = data_d1[103:96];
        7'd14: vec_data_111 = data_d1[111:104];
        7'd15: vec_data_111 = data_d1[119:112];
        7'd16: vec_data_111 = data_d1[127:120];
        7'd17: vec_data_111 = data_d1[135:128];
        7'd18: vec_data_111 = data_d1[143:136];
        7'd19: vec_data_111 = data_d1[151:144];
        7'd20: vec_data_111 = data_d1[159:152];
        7'd21: vec_data_111 = data_d1[167:160];
        7'd22: vec_data_111 = data_d1[175:168];
        7'd23: vec_data_111 = data_d1[183:176];
        7'd24: vec_data_111 = data_d1[191:184];
        7'd25: vec_data_111 = data_d1[199:192];
        7'd26: vec_data_111 = data_d1[207:200];
        7'd27: vec_data_111 = data_d1[215:208];
        7'd28: vec_data_111 = data_d1[223:216];
        7'd29: vec_data_111 = data_d1[231:224];
        7'd30: vec_data_111 = data_d1[239:232];
        7'd31: vec_data_111 = data_d1[247:240];
        7'd32: vec_data_111 = data_d1[255:248];
        7'd33: vec_data_111 = data_d1[263:256];
        7'd34: vec_data_111 = data_d1[271:264];
        7'd35: vec_data_111 = data_d1[279:272];
        7'd36: vec_data_111 = data_d1[287:280];
        7'd37: vec_data_111 = data_d1[295:288];
        7'd38: vec_data_111 = data_d1[303:296];
        7'd39: vec_data_111 = data_d1[311:304];
        7'd40: vec_data_111 = data_d1[319:312];
        7'd41: vec_data_111 = data_d1[327:320];
        7'd42: vec_data_111 = data_d1[335:328];
        7'd43: vec_data_111 = data_d1[343:336];
        7'd44: vec_data_111 = data_d1[351:344];
        7'd45: vec_data_111 = data_d1[359:352];
        7'd46: vec_data_111 = data_d1[367:360];
        7'd47: vec_data_111 = data_d1[375:368];
        7'd48: vec_data_111 = data_d1[383:376];
        7'd49: vec_data_111 = data_d1[391:384];
        7'd50: vec_data_111 = data_d1[399:392];
        7'd51: vec_data_111 = data_d1[407:400];
        7'd52: vec_data_111 = data_d1[415:408];
        7'd53: vec_data_111 = data_d1[423:416];
        7'd54: vec_data_111 = data_d1[431:424];
        7'd55: vec_data_111 = data_d1[439:432];
        7'd56: vec_data_111 = data_d1[447:440];
        7'd57: vec_data_111 = data_d1[455:448];
        7'd58: vec_data_111 = data_d1[463:456];
        7'd59: vec_data_111 = data_d1[471:464];
        7'd60: vec_data_111 = data_d1[479:472];
        7'd61: vec_data_111 = data_d1[487:480];
        7'd62: vec_data_111 = data_d1[495:488];
        7'd63: vec_data_111 = data_d1[503:496];
        7'd64: vec_data_111 = data_d1[511:504];
        7'd65: vec_data_111 = data_d1[519:512];
        7'd66: vec_data_111 = data_d1[527:520];
        7'd67: vec_data_111 = data_d1[535:528];
        7'd68: vec_data_111 = data_d1[543:536];
        7'd69: vec_data_111 = data_d1[551:544];
        7'd70: vec_data_111 = data_d1[559:552];
        7'd71: vec_data_111 = data_d1[567:560];
        7'd72: vec_data_111 = data_d1[575:568];
        7'd73: vec_data_111 = data_d1[583:576];
        7'd74: vec_data_111 = data_d1[591:584];
        7'd75: vec_data_111 = data_d1[599:592];
        7'd76: vec_data_111 = data_d1[607:600];
        7'd77: vec_data_111 = data_d1[615:608];
        7'd78: vec_data_111 = data_d1[623:616];
        7'd79: vec_data_111 = data_d1[631:624];
        7'd80: vec_data_111 = data_d1[639:632];
        7'd81: vec_data_111 = data_d1[647:640];
        7'd82: vec_data_111 = data_d1[655:648];
        7'd83: vec_data_111 = data_d1[663:656];
        7'd84: vec_data_111 = data_d1[671:664];
        7'd85: vec_data_111 = data_d1[679:672];
        7'd86: vec_data_111 = data_d1[687:680];
        7'd87: vec_data_111 = data_d1[695:688];
        7'd88: vec_data_111 = data_d1[703:696];
        7'd89: vec_data_111 = data_d1[711:704];
        7'd90: vec_data_111 = data_d1[719:712];
        7'd91: vec_data_111 = data_d1[727:720];
        7'd92: vec_data_111 = data_d1[735:728];
        7'd93: vec_data_111 = data_d1[743:736];
        7'd94: vec_data_111 = data_d1[751:744];
        7'd95: vec_data_111 = data_d1[759:752];
        7'd96: vec_data_111 = data_d1[767:760];
        7'd97: vec_data_111 = data_d1[775:768];
        7'd98: vec_data_111 = data_d1[783:776];
        7'd99: vec_data_111 = data_d1[791:784];
        7'd100: vec_data_111 = data_d1[799:792];
        7'd101: vec_data_111 = data_d1[807:800];
        7'd102: vec_data_111 = data_d1[815:808];
        7'd103: vec_data_111 = data_d1[823:816];
        7'd104: vec_data_111 = data_d1[831:824];
        7'd105: vec_data_111 = data_d1[839:832];
        7'd106: vec_data_111 = data_d1[847:840];
        7'd107: vec_data_111 = data_d1[855:848];
        7'd108: vec_data_111 = data_d1[863:856];
        7'd109: vec_data_111 = data_d1[871:864];
        7'd110: vec_data_111 = data_d1[879:872];
        7'd111: vec_data_111 = data_d1[887:880];
        7'd112: vec_data_111 = data_d1[895:888];
    endcase
end

always @(
  vec_sum_112_d1
  or data_d1
  ) begin
    vec_data_112 = 8'b0;
    case(vec_sum_112_d1)
        7'd1: vec_data_112 = data_d1[7:0];
        7'd2: vec_data_112 = data_d1[15:8];
        7'd3: vec_data_112 = data_d1[23:16];
        7'd4: vec_data_112 = data_d1[31:24];
        7'd5: vec_data_112 = data_d1[39:32];
        7'd6: vec_data_112 = data_d1[47:40];
        7'd7: vec_data_112 = data_d1[55:48];
        7'd8: vec_data_112 = data_d1[63:56];
        7'd9: vec_data_112 = data_d1[71:64];
        7'd10: vec_data_112 = data_d1[79:72];
        7'd11: vec_data_112 = data_d1[87:80];
        7'd12: vec_data_112 = data_d1[95:88];
        7'd13: vec_data_112 = data_d1[103:96];
        7'd14: vec_data_112 = data_d1[111:104];
        7'd15: vec_data_112 = data_d1[119:112];
        7'd16: vec_data_112 = data_d1[127:120];
        7'd17: vec_data_112 = data_d1[135:128];
        7'd18: vec_data_112 = data_d1[143:136];
        7'd19: vec_data_112 = data_d1[151:144];
        7'd20: vec_data_112 = data_d1[159:152];
        7'd21: vec_data_112 = data_d1[167:160];
        7'd22: vec_data_112 = data_d1[175:168];
        7'd23: vec_data_112 = data_d1[183:176];
        7'd24: vec_data_112 = data_d1[191:184];
        7'd25: vec_data_112 = data_d1[199:192];
        7'd26: vec_data_112 = data_d1[207:200];
        7'd27: vec_data_112 = data_d1[215:208];
        7'd28: vec_data_112 = data_d1[223:216];
        7'd29: vec_data_112 = data_d1[231:224];
        7'd30: vec_data_112 = data_d1[239:232];
        7'd31: vec_data_112 = data_d1[247:240];
        7'd32: vec_data_112 = data_d1[255:248];
        7'd33: vec_data_112 = data_d1[263:256];
        7'd34: vec_data_112 = data_d1[271:264];
        7'd35: vec_data_112 = data_d1[279:272];
        7'd36: vec_data_112 = data_d1[287:280];
        7'd37: vec_data_112 = data_d1[295:288];
        7'd38: vec_data_112 = data_d1[303:296];
        7'd39: vec_data_112 = data_d1[311:304];
        7'd40: vec_data_112 = data_d1[319:312];
        7'd41: vec_data_112 = data_d1[327:320];
        7'd42: vec_data_112 = data_d1[335:328];
        7'd43: vec_data_112 = data_d1[343:336];
        7'd44: vec_data_112 = data_d1[351:344];
        7'd45: vec_data_112 = data_d1[359:352];
        7'd46: vec_data_112 = data_d1[367:360];
        7'd47: vec_data_112 = data_d1[375:368];
        7'd48: vec_data_112 = data_d1[383:376];
        7'd49: vec_data_112 = data_d1[391:384];
        7'd50: vec_data_112 = data_d1[399:392];
        7'd51: vec_data_112 = data_d1[407:400];
        7'd52: vec_data_112 = data_d1[415:408];
        7'd53: vec_data_112 = data_d1[423:416];
        7'd54: vec_data_112 = data_d1[431:424];
        7'd55: vec_data_112 = data_d1[439:432];
        7'd56: vec_data_112 = data_d1[447:440];
        7'd57: vec_data_112 = data_d1[455:448];
        7'd58: vec_data_112 = data_d1[463:456];
        7'd59: vec_data_112 = data_d1[471:464];
        7'd60: vec_data_112 = data_d1[479:472];
        7'd61: vec_data_112 = data_d1[487:480];
        7'd62: vec_data_112 = data_d1[495:488];
        7'd63: vec_data_112 = data_d1[503:496];
        7'd64: vec_data_112 = data_d1[511:504];
        7'd65: vec_data_112 = data_d1[519:512];
        7'd66: vec_data_112 = data_d1[527:520];
        7'd67: vec_data_112 = data_d1[535:528];
        7'd68: vec_data_112 = data_d1[543:536];
        7'd69: vec_data_112 = data_d1[551:544];
        7'd70: vec_data_112 = data_d1[559:552];
        7'd71: vec_data_112 = data_d1[567:560];
        7'd72: vec_data_112 = data_d1[575:568];
        7'd73: vec_data_112 = data_d1[583:576];
        7'd74: vec_data_112 = data_d1[591:584];
        7'd75: vec_data_112 = data_d1[599:592];
        7'd76: vec_data_112 = data_d1[607:600];
        7'd77: vec_data_112 = data_d1[615:608];
        7'd78: vec_data_112 = data_d1[623:616];
        7'd79: vec_data_112 = data_d1[631:624];
        7'd80: vec_data_112 = data_d1[639:632];
        7'd81: vec_data_112 = data_d1[647:640];
        7'd82: vec_data_112 = data_d1[655:648];
        7'd83: vec_data_112 = data_d1[663:656];
        7'd84: vec_data_112 = data_d1[671:664];
        7'd85: vec_data_112 = data_d1[679:672];
        7'd86: vec_data_112 = data_d1[687:680];
        7'd87: vec_data_112 = data_d1[695:688];
        7'd88: vec_data_112 = data_d1[703:696];
        7'd89: vec_data_112 = data_d1[711:704];
        7'd90: vec_data_112 = data_d1[719:712];
        7'd91: vec_data_112 = data_d1[727:720];
        7'd92: vec_data_112 = data_d1[735:728];
        7'd93: vec_data_112 = data_d1[743:736];
        7'd94: vec_data_112 = data_d1[751:744];
        7'd95: vec_data_112 = data_d1[759:752];
        7'd96: vec_data_112 = data_d1[767:760];
        7'd97: vec_data_112 = data_d1[775:768];
        7'd98: vec_data_112 = data_d1[783:776];
        7'd99: vec_data_112 = data_d1[791:784];
        7'd100: vec_data_112 = data_d1[799:792];
        7'd101: vec_data_112 = data_d1[807:800];
        7'd102: vec_data_112 = data_d1[815:808];
        7'd103: vec_data_112 = data_d1[823:816];
        7'd104: vec_data_112 = data_d1[831:824];
        7'd105: vec_data_112 = data_d1[839:832];
        7'd106: vec_data_112 = data_d1[847:840];
        7'd107: vec_data_112 = data_d1[855:848];
        7'd108: vec_data_112 = data_d1[863:856];
        7'd109: vec_data_112 = data_d1[871:864];
        7'd110: vec_data_112 = data_d1[879:872];
        7'd111: vec_data_112 = data_d1[887:880];
        7'd112: vec_data_112 = data_d1[895:888];
        7'd113: vec_data_112 = data_d1[903:896];
    endcase
end

always @(
  vec_sum_113_d1
  or data_d1
  ) begin
    vec_data_113 = 8'b0;
    case(vec_sum_113_d1)
        7'd1: vec_data_113 = data_d1[7:0];
        7'd2: vec_data_113 = data_d1[15:8];
        7'd3: vec_data_113 = data_d1[23:16];
        7'd4: vec_data_113 = data_d1[31:24];
        7'd5: vec_data_113 = data_d1[39:32];
        7'd6: vec_data_113 = data_d1[47:40];
        7'd7: vec_data_113 = data_d1[55:48];
        7'd8: vec_data_113 = data_d1[63:56];
        7'd9: vec_data_113 = data_d1[71:64];
        7'd10: vec_data_113 = data_d1[79:72];
        7'd11: vec_data_113 = data_d1[87:80];
        7'd12: vec_data_113 = data_d1[95:88];
        7'd13: vec_data_113 = data_d1[103:96];
        7'd14: vec_data_113 = data_d1[111:104];
        7'd15: vec_data_113 = data_d1[119:112];
        7'd16: vec_data_113 = data_d1[127:120];
        7'd17: vec_data_113 = data_d1[135:128];
        7'd18: vec_data_113 = data_d1[143:136];
        7'd19: vec_data_113 = data_d1[151:144];
        7'd20: vec_data_113 = data_d1[159:152];
        7'd21: vec_data_113 = data_d1[167:160];
        7'd22: vec_data_113 = data_d1[175:168];
        7'd23: vec_data_113 = data_d1[183:176];
        7'd24: vec_data_113 = data_d1[191:184];
        7'd25: vec_data_113 = data_d1[199:192];
        7'd26: vec_data_113 = data_d1[207:200];
        7'd27: vec_data_113 = data_d1[215:208];
        7'd28: vec_data_113 = data_d1[223:216];
        7'd29: vec_data_113 = data_d1[231:224];
        7'd30: vec_data_113 = data_d1[239:232];
        7'd31: vec_data_113 = data_d1[247:240];
        7'd32: vec_data_113 = data_d1[255:248];
        7'd33: vec_data_113 = data_d1[263:256];
        7'd34: vec_data_113 = data_d1[271:264];
        7'd35: vec_data_113 = data_d1[279:272];
        7'd36: vec_data_113 = data_d1[287:280];
        7'd37: vec_data_113 = data_d1[295:288];
        7'd38: vec_data_113 = data_d1[303:296];
        7'd39: vec_data_113 = data_d1[311:304];
        7'd40: vec_data_113 = data_d1[319:312];
        7'd41: vec_data_113 = data_d1[327:320];
        7'd42: vec_data_113 = data_d1[335:328];
        7'd43: vec_data_113 = data_d1[343:336];
        7'd44: vec_data_113 = data_d1[351:344];
        7'd45: vec_data_113 = data_d1[359:352];
        7'd46: vec_data_113 = data_d1[367:360];
        7'd47: vec_data_113 = data_d1[375:368];
        7'd48: vec_data_113 = data_d1[383:376];
        7'd49: vec_data_113 = data_d1[391:384];
        7'd50: vec_data_113 = data_d1[399:392];
        7'd51: vec_data_113 = data_d1[407:400];
        7'd52: vec_data_113 = data_d1[415:408];
        7'd53: vec_data_113 = data_d1[423:416];
        7'd54: vec_data_113 = data_d1[431:424];
        7'd55: vec_data_113 = data_d1[439:432];
        7'd56: vec_data_113 = data_d1[447:440];
        7'd57: vec_data_113 = data_d1[455:448];
        7'd58: vec_data_113 = data_d1[463:456];
        7'd59: vec_data_113 = data_d1[471:464];
        7'd60: vec_data_113 = data_d1[479:472];
        7'd61: vec_data_113 = data_d1[487:480];
        7'd62: vec_data_113 = data_d1[495:488];
        7'd63: vec_data_113 = data_d1[503:496];
        7'd64: vec_data_113 = data_d1[511:504];
        7'd65: vec_data_113 = data_d1[519:512];
        7'd66: vec_data_113 = data_d1[527:520];
        7'd67: vec_data_113 = data_d1[535:528];
        7'd68: vec_data_113 = data_d1[543:536];
        7'd69: vec_data_113 = data_d1[551:544];
        7'd70: vec_data_113 = data_d1[559:552];
        7'd71: vec_data_113 = data_d1[567:560];
        7'd72: vec_data_113 = data_d1[575:568];
        7'd73: vec_data_113 = data_d1[583:576];
        7'd74: vec_data_113 = data_d1[591:584];
        7'd75: vec_data_113 = data_d1[599:592];
        7'd76: vec_data_113 = data_d1[607:600];
        7'd77: vec_data_113 = data_d1[615:608];
        7'd78: vec_data_113 = data_d1[623:616];
        7'd79: vec_data_113 = data_d1[631:624];
        7'd80: vec_data_113 = data_d1[639:632];
        7'd81: vec_data_113 = data_d1[647:640];
        7'd82: vec_data_113 = data_d1[655:648];
        7'd83: vec_data_113 = data_d1[663:656];
        7'd84: vec_data_113 = data_d1[671:664];
        7'd85: vec_data_113 = data_d1[679:672];
        7'd86: vec_data_113 = data_d1[687:680];
        7'd87: vec_data_113 = data_d1[695:688];
        7'd88: vec_data_113 = data_d1[703:696];
        7'd89: vec_data_113 = data_d1[711:704];
        7'd90: vec_data_113 = data_d1[719:712];
        7'd91: vec_data_113 = data_d1[727:720];
        7'd92: vec_data_113 = data_d1[735:728];
        7'd93: vec_data_113 = data_d1[743:736];
        7'd94: vec_data_113 = data_d1[751:744];
        7'd95: vec_data_113 = data_d1[759:752];
        7'd96: vec_data_113 = data_d1[767:760];
        7'd97: vec_data_113 = data_d1[775:768];
        7'd98: vec_data_113 = data_d1[783:776];
        7'd99: vec_data_113 = data_d1[791:784];
        7'd100: vec_data_113 = data_d1[799:792];
        7'd101: vec_data_113 = data_d1[807:800];
        7'd102: vec_data_113 = data_d1[815:808];
        7'd103: vec_data_113 = data_d1[823:816];
        7'd104: vec_data_113 = data_d1[831:824];
        7'd105: vec_data_113 = data_d1[839:832];
        7'd106: vec_data_113 = data_d1[847:840];
        7'd107: vec_data_113 = data_d1[855:848];
        7'd108: vec_data_113 = data_d1[863:856];
        7'd109: vec_data_113 = data_d1[871:864];
        7'd110: vec_data_113 = data_d1[879:872];
        7'd111: vec_data_113 = data_d1[887:880];
        7'd112: vec_data_113 = data_d1[895:888];
        7'd113: vec_data_113 = data_d1[903:896];
        7'd114: vec_data_113 = data_d1[911:904];
    endcase
end

always @(
  vec_sum_114_d1
  or data_d1
  ) begin
    vec_data_114 = 8'b0;
    case(vec_sum_114_d1)
        7'd1: vec_data_114 = data_d1[7:0];
        7'd2: vec_data_114 = data_d1[15:8];
        7'd3: vec_data_114 = data_d1[23:16];
        7'd4: vec_data_114 = data_d1[31:24];
        7'd5: vec_data_114 = data_d1[39:32];
        7'd6: vec_data_114 = data_d1[47:40];
        7'd7: vec_data_114 = data_d1[55:48];
        7'd8: vec_data_114 = data_d1[63:56];
        7'd9: vec_data_114 = data_d1[71:64];
        7'd10: vec_data_114 = data_d1[79:72];
        7'd11: vec_data_114 = data_d1[87:80];
        7'd12: vec_data_114 = data_d1[95:88];
        7'd13: vec_data_114 = data_d1[103:96];
        7'd14: vec_data_114 = data_d1[111:104];
        7'd15: vec_data_114 = data_d1[119:112];
        7'd16: vec_data_114 = data_d1[127:120];
        7'd17: vec_data_114 = data_d1[135:128];
        7'd18: vec_data_114 = data_d1[143:136];
        7'd19: vec_data_114 = data_d1[151:144];
        7'd20: vec_data_114 = data_d1[159:152];
        7'd21: vec_data_114 = data_d1[167:160];
        7'd22: vec_data_114 = data_d1[175:168];
        7'd23: vec_data_114 = data_d1[183:176];
        7'd24: vec_data_114 = data_d1[191:184];
        7'd25: vec_data_114 = data_d1[199:192];
        7'd26: vec_data_114 = data_d1[207:200];
        7'd27: vec_data_114 = data_d1[215:208];
        7'd28: vec_data_114 = data_d1[223:216];
        7'd29: vec_data_114 = data_d1[231:224];
        7'd30: vec_data_114 = data_d1[239:232];
        7'd31: vec_data_114 = data_d1[247:240];
        7'd32: vec_data_114 = data_d1[255:248];
        7'd33: vec_data_114 = data_d1[263:256];
        7'd34: vec_data_114 = data_d1[271:264];
        7'd35: vec_data_114 = data_d1[279:272];
        7'd36: vec_data_114 = data_d1[287:280];
        7'd37: vec_data_114 = data_d1[295:288];
        7'd38: vec_data_114 = data_d1[303:296];
        7'd39: vec_data_114 = data_d1[311:304];
        7'd40: vec_data_114 = data_d1[319:312];
        7'd41: vec_data_114 = data_d1[327:320];
        7'd42: vec_data_114 = data_d1[335:328];
        7'd43: vec_data_114 = data_d1[343:336];
        7'd44: vec_data_114 = data_d1[351:344];
        7'd45: vec_data_114 = data_d1[359:352];
        7'd46: vec_data_114 = data_d1[367:360];
        7'd47: vec_data_114 = data_d1[375:368];
        7'd48: vec_data_114 = data_d1[383:376];
        7'd49: vec_data_114 = data_d1[391:384];
        7'd50: vec_data_114 = data_d1[399:392];
        7'd51: vec_data_114 = data_d1[407:400];
        7'd52: vec_data_114 = data_d1[415:408];
        7'd53: vec_data_114 = data_d1[423:416];
        7'd54: vec_data_114 = data_d1[431:424];
        7'd55: vec_data_114 = data_d1[439:432];
        7'd56: vec_data_114 = data_d1[447:440];
        7'd57: vec_data_114 = data_d1[455:448];
        7'd58: vec_data_114 = data_d1[463:456];
        7'd59: vec_data_114 = data_d1[471:464];
        7'd60: vec_data_114 = data_d1[479:472];
        7'd61: vec_data_114 = data_d1[487:480];
        7'd62: vec_data_114 = data_d1[495:488];
        7'd63: vec_data_114 = data_d1[503:496];
        7'd64: vec_data_114 = data_d1[511:504];
        7'd65: vec_data_114 = data_d1[519:512];
        7'd66: vec_data_114 = data_d1[527:520];
        7'd67: vec_data_114 = data_d1[535:528];
        7'd68: vec_data_114 = data_d1[543:536];
        7'd69: vec_data_114 = data_d1[551:544];
        7'd70: vec_data_114 = data_d1[559:552];
        7'd71: vec_data_114 = data_d1[567:560];
        7'd72: vec_data_114 = data_d1[575:568];
        7'd73: vec_data_114 = data_d1[583:576];
        7'd74: vec_data_114 = data_d1[591:584];
        7'd75: vec_data_114 = data_d1[599:592];
        7'd76: vec_data_114 = data_d1[607:600];
        7'd77: vec_data_114 = data_d1[615:608];
        7'd78: vec_data_114 = data_d1[623:616];
        7'd79: vec_data_114 = data_d1[631:624];
        7'd80: vec_data_114 = data_d1[639:632];
        7'd81: vec_data_114 = data_d1[647:640];
        7'd82: vec_data_114 = data_d1[655:648];
        7'd83: vec_data_114 = data_d1[663:656];
        7'd84: vec_data_114 = data_d1[671:664];
        7'd85: vec_data_114 = data_d1[679:672];
        7'd86: vec_data_114 = data_d1[687:680];
        7'd87: vec_data_114 = data_d1[695:688];
        7'd88: vec_data_114 = data_d1[703:696];
        7'd89: vec_data_114 = data_d1[711:704];
        7'd90: vec_data_114 = data_d1[719:712];
        7'd91: vec_data_114 = data_d1[727:720];
        7'd92: vec_data_114 = data_d1[735:728];
        7'd93: vec_data_114 = data_d1[743:736];
        7'd94: vec_data_114 = data_d1[751:744];
        7'd95: vec_data_114 = data_d1[759:752];
        7'd96: vec_data_114 = data_d1[767:760];
        7'd97: vec_data_114 = data_d1[775:768];
        7'd98: vec_data_114 = data_d1[783:776];
        7'd99: vec_data_114 = data_d1[791:784];
        7'd100: vec_data_114 = data_d1[799:792];
        7'd101: vec_data_114 = data_d1[807:800];
        7'd102: vec_data_114 = data_d1[815:808];
        7'd103: vec_data_114 = data_d1[823:816];
        7'd104: vec_data_114 = data_d1[831:824];
        7'd105: vec_data_114 = data_d1[839:832];
        7'd106: vec_data_114 = data_d1[847:840];
        7'd107: vec_data_114 = data_d1[855:848];
        7'd108: vec_data_114 = data_d1[863:856];
        7'd109: vec_data_114 = data_d1[871:864];
        7'd110: vec_data_114 = data_d1[879:872];
        7'd111: vec_data_114 = data_d1[887:880];
        7'd112: vec_data_114 = data_d1[895:888];
        7'd113: vec_data_114 = data_d1[903:896];
        7'd114: vec_data_114 = data_d1[911:904];
        7'd115: vec_data_114 = data_d1[919:912];
    endcase
end

always @(
  vec_sum_115_d1
  or data_d1
  ) begin
    vec_data_115 = 8'b0;
    case(vec_sum_115_d1)
        7'd1: vec_data_115 = data_d1[7:0];
        7'd2: vec_data_115 = data_d1[15:8];
        7'd3: vec_data_115 = data_d1[23:16];
        7'd4: vec_data_115 = data_d1[31:24];
        7'd5: vec_data_115 = data_d1[39:32];
        7'd6: vec_data_115 = data_d1[47:40];
        7'd7: vec_data_115 = data_d1[55:48];
        7'd8: vec_data_115 = data_d1[63:56];
        7'd9: vec_data_115 = data_d1[71:64];
        7'd10: vec_data_115 = data_d1[79:72];
        7'd11: vec_data_115 = data_d1[87:80];
        7'd12: vec_data_115 = data_d1[95:88];
        7'd13: vec_data_115 = data_d1[103:96];
        7'd14: vec_data_115 = data_d1[111:104];
        7'd15: vec_data_115 = data_d1[119:112];
        7'd16: vec_data_115 = data_d1[127:120];
        7'd17: vec_data_115 = data_d1[135:128];
        7'd18: vec_data_115 = data_d1[143:136];
        7'd19: vec_data_115 = data_d1[151:144];
        7'd20: vec_data_115 = data_d1[159:152];
        7'd21: vec_data_115 = data_d1[167:160];
        7'd22: vec_data_115 = data_d1[175:168];
        7'd23: vec_data_115 = data_d1[183:176];
        7'd24: vec_data_115 = data_d1[191:184];
        7'd25: vec_data_115 = data_d1[199:192];
        7'd26: vec_data_115 = data_d1[207:200];
        7'd27: vec_data_115 = data_d1[215:208];
        7'd28: vec_data_115 = data_d1[223:216];
        7'd29: vec_data_115 = data_d1[231:224];
        7'd30: vec_data_115 = data_d1[239:232];
        7'd31: vec_data_115 = data_d1[247:240];
        7'd32: vec_data_115 = data_d1[255:248];
        7'd33: vec_data_115 = data_d1[263:256];
        7'd34: vec_data_115 = data_d1[271:264];
        7'd35: vec_data_115 = data_d1[279:272];
        7'd36: vec_data_115 = data_d1[287:280];
        7'd37: vec_data_115 = data_d1[295:288];
        7'd38: vec_data_115 = data_d1[303:296];
        7'd39: vec_data_115 = data_d1[311:304];
        7'd40: vec_data_115 = data_d1[319:312];
        7'd41: vec_data_115 = data_d1[327:320];
        7'd42: vec_data_115 = data_d1[335:328];
        7'd43: vec_data_115 = data_d1[343:336];
        7'd44: vec_data_115 = data_d1[351:344];
        7'd45: vec_data_115 = data_d1[359:352];
        7'd46: vec_data_115 = data_d1[367:360];
        7'd47: vec_data_115 = data_d1[375:368];
        7'd48: vec_data_115 = data_d1[383:376];
        7'd49: vec_data_115 = data_d1[391:384];
        7'd50: vec_data_115 = data_d1[399:392];
        7'd51: vec_data_115 = data_d1[407:400];
        7'd52: vec_data_115 = data_d1[415:408];
        7'd53: vec_data_115 = data_d1[423:416];
        7'd54: vec_data_115 = data_d1[431:424];
        7'd55: vec_data_115 = data_d1[439:432];
        7'd56: vec_data_115 = data_d1[447:440];
        7'd57: vec_data_115 = data_d1[455:448];
        7'd58: vec_data_115 = data_d1[463:456];
        7'd59: vec_data_115 = data_d1[471:464];
        7'd60: vec_data_115 = data_d1[479:472];
        7'd61: vec_data_115 = data_d1[487:480];
        7'd62: vec_data_115 = data_d1[495:488];
        7'd63: vec_data_115 = data_d1[503:496];
        7'd64: vec_data_115 = data_d1[511:504];
        7'd65: vec_data_115 = data_d1[519:512];
        7'd66: vec_data_115 = data_d1[527:520];
        7'd67: vec_data_115 = data_d1[535:528];
        7'd68: vec_data_115 = data_d1[543:536];
        7'd69: vec_data_115 = data_d1[551:544];
        7'd70: vec_data_115 = data_d1[559:552];
        7'd71: vec_data_115 = data_d1[567:560];
        7'd72: vec_data_115 = data_d1[575:568];
        7'd73: vec_data_115 = data_d1[583:576];
        7'd74: vec_data_115 = data_d1[591:584];
        7'd75: vec_data_115 = data_d1[599:592];
        7'd76: vec_data_115 = data_d1[607:600];
        7'd77: vec_data_115 = data_d1[615:608];
        7'd78: vec_data_115 = data_d1[623:616];
        7'd79: vec_data_115 = data_d1[631:624];
        7'd80: vec_data_115 = data_d1[639:632];
        7'd81: vec_data_115 = data_d1[647:640];
        7'd82: vec_data_115 = data_d1[655:648];
        7'd83: vec_data_115 = data_d1[663:656];
        7'd84: vec_data_115 = data_d1[671:664];
        7'd85: vec_data_115 = data_d1[679:672];
        7'd86: vec_data_115 = data_d1[687:680];
        7'd87: vec_data_115 = data_d1[695:688];
        7'd88: vec_data_115 = data_d1[703:696];
        7'd89: vec_data_115 = data_d1[711:704];
        7'd90: vec_data_115 = data_d1[719:712];
        7'd91: vec_data_115 = data_d1[727:720];
        7'd92: vec_data_115 = data_d1[735:728];
        7'd93: vec_data_115 = data_d1[743:736];
        7'd94: vec_data_115 = data_d1[751:744];
        7'd95: vec_data_115 = data_d1[759:752];
        7'd96: vec_data_115 = data_d1[767:760];
        7'd97: vec_data_115 = data_d1[775:768];
        7'd98: vec_data_115 = data_d1[783:776];
        7'd99: vec_data_115 = data_d1[791:784];
        7'd100: vec_data_115 = data_d1[799:792];
        7'd101: vec_data_115 = data_d1[807:800];
        7'd102: vec_data_115 = data_d1[815:808];
        7'd103: vec_data_115 = data_d1[823:816];
        7'd104: vec_data_115 = data_d1[831:824];
        7'd105: vec_data_115 = data_d1[839:832];
        7'd106: vec_data_115 = data_d1[847:840];
        7'd107: vec_data_115 = data_d1[855:848];
        7'd108: vec_data_115 = data_d1[863:856];
        7'd109: vec_data_115 = data_d1[871:864];
        7'd110: vec_data_115 = data_d1[879:872];
        7'd111: vec_data_115 = data_d1[887:880];
        7'd112: vec_data_115 = data_d1[895:888];
        7'd113: vec_data_115 = data_d1[903:896];
        7'd114: vec_data_115 = data_d1[911:904];
        7'd115: vec_data_115 = data_d1[919:912];
        7'd116: vec_data_115 = data_d1[927:920];
    endcase
end

always @(
  vec_sum_116_d1
  or data_d1
  ) begin
    vec_data_116 = 8'b0;
    case(vec_sum_116_d1)
        7'd1: vec_data_116 = data_d1[7:0];
        7'd2: vec_data_116 = data_d1[15:8];
        7'd3: vec_data_116 = data_d1[23:16];
        7'd4: vec_data_116 = data_d1[31:24];
        7'd5: vec_data_116 = data_d1[39:32];
        7'd6: vec_data_116 = data_d1[47:40];
        7'd7: vec_data_116 = data_d1[55:48];
        7'd8: vec_data_116 = data_d1[63:56];
        7'd9: vec_data_116 = data_d1[71:64];
        7'd10: vec_data_116 = data_d1[79:72];
        7'd11: vec_data_116 = data_d1[87:80];
        7'd12: vec_data_116 = data_d1[95:88];
        7'd13: vec_data_116 = data_d1[103:96];
        7'd14: vec_data_116 = data_d1[111:104];
        7'd15: vec_data_116 = data_d1[119:112];
        7'd16: vec_data_116 = data_d1[127:120];
        7'd17: vec_data_116 = data_d1[135:128];
        7'd18: vec_data_116 = data_d1[143:136];
        7'd19: vec_data_116 = data_d1[151:144];
        7'd20: vec_data_116 = data_d1[159:152];
        7'd21: vec_data_116 = data_d1[167:160];
        7'd22: vec_data_116 = data_d1[175:168];
        7'd23: vec_data_116 = data_d1[183:176];
        7'd24: vec_data_116 = data_d1[191:184];
        7'd25: vec_data_116 = data_d1[199:192];
        7'd26: vec_data_116 = data_d1[207:200];
        7'd27: vec_data_116 = data_d1[215:208];
        7'd28: vec_data_116 = data_d1[223:216];
        7'd29: vec_data_116 = data_d1[231:224];
        7'd30: vec_data_116 = data_d1[239:232];
        7'd31: vec_data_116 = data_d1[247:240];
        7'd32: vec_data_116 = data_d1[255:248];
        7'd33: vec_data_116 = data_d1[263:256];
        7'd34: vec_data_116 = data_d1[271:264];
        7'd35: vec_data_116 = data_d1[279:272];
        7'd36: vec_data_116 = data_d1[287:280];
        7'd37: vec_data_116 = data_d1[295:288];
        7'd38: vec_data_116 = data_d1[303:296];
        7'd39: vec_data_116 = data_d1[311:304];
        7'd40: vec_data_116 = data_d1[319:312];
        7'd41: vec_data_116 = data_d1[327:320];
        7'd42: vec_data_116 = data_d1[335:328];
        7'd43: vec_data_116 = data_d1[343:336];
        7'd44: vec_data_116 = data_d1[351:344];
        7'd45: vec_data_116 = data_d1[359:352];
        7'd46: vec_data_116 = data_d1[367:360];
        7'd47: vec_data_116 = data_d1[375:368];
        7'd48: vec_data_116 = data_d1[383:376];
        7'd49: vec_data_116 = data_d1[391:384];
        7'd50: vec_data_116 = data_d1[399:392];
        7'd51: vec_data_116 = data_d1[407:400];
        7'd52: vec_data_116 = data_d1[415:408];
        7'd53: vec_data_116 = data_d1[423:416];
        7'd54: vec_data_116 = data_d1[431:424];
        7'd55: vec_data_116 = data_d1[439:432];
        7'd56: vec_data_116 = data_d1[447:440];
        7'd57: vec_data_116 = data_d1[455:448];
        7'd58: vec_data_116 = data_d1[463:456];
        7'd59: vec_data_116 = data_d1[471:464];
        7'd60: vec_data_116 = data_d1[479:472];
        7'd61: vec_data_116 = data_d1[487:480];
        7'd62: vec_data_116 = data_d1[495:488];
        7'd63: vec_data_116 = data_d1[503:496];
        7'd64: vec_data_116 = data_d1[511:504];
        7'd65: vec_data_116 = data_d1[519:512];
        7'd66: vec_data_116 = data_d1[527:520];
        7'd67: vec_data_116 = data_d1[535:528];
        7'd68: vec_data_116 = data_d1[543:536];
        7'd69: vec_data_116 = data_d1[551:544];
        7'd70: vec_data_116 = data_d1[559:552];
        7'd71: vec_data_116 = data_d1[567:560];
        7'd72: vec_data_116 = data_d1[575:568];
        7'd73: vec_data_116 = data_d1[583:576];
        7'd74: vec_data_116 = data_d1[591:584];
        7'd75: vec_data_116 = data_d1[599:592];
        7'd76: vec_data_116 = data_d1[607:600];
        7'd77: vec_data_116 = data_d1[615:608];
        7'd78: vec_data_116 = data_d1[623:616];
        7'd79: vec_data_116 = data_d1[631:624];
        7'd80: vec_data_116 = data_d1[639:632];
        7'd81: vec_data_116 = data_d1[647:640];
        7'd82: vec_data_116 = data_d1[655:648];
        7'd83: vec_data_116 = data_d1[663:656];
        7'd84: vec_data_116 = data_d1[671:664];
        7'd85: vec_data_116 = data_d1[679:672];
        7'd86: vec_data_116 = data_d1[687:680];
        7'd87: vec_data_116 = data_d1[695:688];
        7'd88: vec_data_116 = data_d1[703:696];
        7'd89: vec_data_116 = data_d1[711:704];
        7'd90: vec_data_116 = data_d1[719:712];
        7'd91: vec_data_116 = data_d1[727:720];
        7'd92: vec_data_116 = data_d1[735:728];
        7'd93: vec_data_116 = data_d1[743:736];
        7'd94: vec_data_116 = data_d1[751:744];
        7'd95: vec_data_116 = data_d1[759:752];
        7'd96: vec_data_116 = data_d1[767:760];
        7'd97: vec_data_116 = data_d1[775:768];
        7'd98: vec_data_116 = data_d1[783:776];
        7'd99: vec_data_116 = data_d1[791:784];
        7'd100: vec_data_116 = data_d1[799:792];
        7'd101: vec_data_116 = data_d1[807:800];
        7'd102: vec_data_116 = data_d1[815:808];
        7'd103: vec_data_116 = data_d1[823:816];
        7'd104: vec_data_116 = data_d1[831:824];
        7'd105: vec_data_116 = data_d1[839:832];
        7'd106: vec_data_116 = data_d1[847:840];
        7'd107: vec_data_116 = data_d1[855:848];
        7'd108: vec_data_116 = data_d1[863:856];
        7'd109: vec_data_116 = data_d1[871:864];
        7'd110: vec_data_116 = data_d1[879:872];
        7'd111: vec_data_116 = data_d1[887:880];
        7'd112: vec_data_116 = data_d1[895:888];
        7'd113: vec_data_116 = data_d1[903:896];
        7'd114: vec_data_116 = data_d1[911:904];
        7'd115: vec_data_116 = data_d1[919:912];
        7'd116: vec_data_116 = data_d1[927:920];
        7'd117: vec_data_116 = data_d1[935:928];
    endcase
end

always @(
  vec_sum_117_d1
  or data_d1
  ) begin
    vec_data_117 = 8'b0;
    case(vec_sum_117_d1)
        7'd1: vec_data_117 = data_d1[7:0];
        7'd2: vec_data_117 = data_d1[15:8];
        7'd3: vec_data_117 = data_d1[23:16];
        7'd4: vec_data_117 = data_d1[31:24];
        7'd5: vec_data_117 = data_d1[39:32];
        7'd6: vec_data_117 = data_d1[47:40];
        7'd7: vec_data_117 = data_d1[55:48];
        7'd8: vec_data_117 = data_d1[63:56];
        7'd9: vec_data_117 = data_d1[71:64];
        7'd10: vec_data_117 = data_d1[79:72];
        7'd11: vec_data_117 = data_d1[87:80];
        7'd12: vec_data_117 = data_d1[95:88];
        7'd13: vec_data_117 = data_d1[103:96];
        7'd14: vec_data_117 = data_d1[111:104];
        7'd15: vec_data_117 = data_d1[119:112];
        7'd16: vec_data_117 = data_d1[127:120];
        7'd17: vec_data_117 = data_d1[135:128];
        7'd18: vec_data_117 = data_d1[143:136];
        7'd19: vec_data_117 = data_d1[151:144];
        7'd20: vec_data_117 = data_d1[159:152];
        7'd21: vec_data_117 = data_d1[167:160];
        7'd22: vec_data_117 = data_d1[175:168];
        7'd23: vec_data_117 = data_d1[183:176];
        7'd24: vec_data_117 = data_d1[191:184];
        7'd25: vec_data_117 = data_d1[199:192];
        7'd26: vec_data_117 = data_d1[207:200];
        7'd27: vec_data_117 = data_d1[215:208];
        7'd28: vec_data_117 = data_d1[223:216];
        7'd29: vec_data_117 = data_d1[231:224];
        7'd30: vec_data_117 = data_d1[239:232];
        7'd31: vec_data_117 = data_d1[247:240];
        7'd32: vec_data_117 = data_d1[255:248];
        7'd33: vec_data_117 = data_d1[263:256];
        7'd34: vec_data_117 = data_d1[271:264];
        7'd35: vec_data_117 = data_d1[279:272];
        7'd36: vec_data_117 = data_d1[287:280];
        7'd37: vec_data_117 = data_d1[295:288];
        7'd38: vec_data_117 = data_d1[303:296];
        7'd39: vec_data_117 = data_d1[311:304];
        7'd40: vec_data_117 = data_d1[319:312];
        7'd41: vec_data_117 = data_d1[327:320];
        7'd42: vec_data_117 = data_d1[335:328];
        7'd43: vec_data_117 = data_d1[343:336];
        7'd44: vec_data_117 = data_d1[351:344];
        7'd45: vec_data_117 = data_d1[359:352];
        7'd46: vec_data_117 = data_d1[367:360];
        7'd47: vec_data_117 = data_d1[375:368];
        7'd48: vec_data_117 = data_d1[383:376];
        7'd49: vec_data_117 = data_d1[391:384];
        7'd50: vec_data_117 = data_d1[399:392];
        7'd51: vec_data_117 = data_d1[407:400];
        7'd52: vec_data_117 = data_d1[415:408];
        7'd53: vec_data_117 = data_d1[423:416];
        7'd54: vec_data_117 = data_d1[431:424];
        7'd55: vec_data_117 = data_d1[439:432];
        7'd56: vec_data_117 = data_d1[447:440];
        7'd57: vec_data_117 = data_d1[455:448];
        7'd58: vec_data_117 = data_d1[463:456];
        7'd59: vec_data_117 = data_d1[471:464];
        7'd60: vec_data_117 = data_d1[479:472];
        7'd61: vec_data_117 = data_d1[487:480];
        7'd62: vec_data_117 = data_d1[495:488];
        7'd63: vec_data_117 = data_d1[503:496];
        7'd64: vec_data_117 = data_d1[511:504];
        7'd65: vec_data_117 = data_d1[519:512];
        7'd66: vec_data_117 = data_d1[527:520];
        7'd67: vec_data_117 = data_d1[535:528];
        7'd68: vec_data_117 = data_d1[543:536];
        7'd69: vec_data_117 = data_d1[551:544];
        7'd70: vec_data_117 = data_d1[559:552];
        7'd71: vec_data_117 = data_d1[567:560];
        7'd72: vec_data_117 = data_d1[575:568];
        7'd73: vec_data_117 = data_d1[583:576];
        7'd74: vec_data_117 = data_d1[591:584];
        7'd75: vec_data_117 = data_d1[599:592];
        7'd76: vec_data_117 = data_d1[607:600];
        7'd77: vec_data_117 = data_d1[615:608];
        7'd78: vec_data_117 = data_d1[623:616];
        7'd79: vec_data_117 = data_d1[631:624];
        7'd80: vec_data_117 = data_d1[639:632];
        7'd81: vec_data_117 = data_d1[647:640];
        7'd82: vec_data_117 = data_d1[655:648];
        7'd83: vec_data_117 = data_d1[663:656];
        7'd84: vec_data_117 = data_d1[671:664];
        7'd85: vec_data_117 = data_d1[679:672];
        7'd86: vec_data_117 = data_d1[687:680];
        7'd87: vec_data_117 = data_d1[695:688];
        7'd88: vec_data_117 = data_d1[703:696];
        7'd89: vec_data_117 = data_d1[711:704];
        7'd90: vec_data_117 = data_d1[719:712];
        7'd91: vec_data_117 = data_d1[727:720];
        7'd92: vec_data_117 = data_d1[735:728];
        7'd93: vec_data_117 = data_d1[743:736];
        7'd94: vec_data_117 = data_d1[751:744];
        7'd95: vec_data_117 = data_d1[759:752];
        7'd96: vec_data_117 = data_d1[767:760];
        7'd97: vec_data_117 = data_d1[775:768];
        7'd98: vec_data_117 = data_d1[783:776];
        7'd99: vec_data_117 = data_d1[791:784];
        7'd100: vec_data_117 = data_d1[799:792];
        7'd101: vec_data_117 = data_d1[807:800];
        7'd102: vec_data_117 = data_d1[815:808];
        7'd103: vec_data_117 = data_d1[823:816];
        7'd104: vec_data_117 = data_d1[831:824];
        7'd105: vec_data_117 = data_d1[839:832];
        7'd106: vec_data_117 = data_d1[847:840];
        7'd107: vec_data_117 = data_d1[855:848];
        7'd108: vec_data_117 = data_d1[863:856];
        7'd109: vec_data_117 = data_d1[871:864];
        7'd110: vec_data_117 = data_d1[879:872];
        7'd111: vec_data_117 = data_d1[887:880];
        7'd112: vec_data_117 = data_d1[895:888];
        7'd113: vec_data_117 = data_d1[903:896];
        7'd114: vec_data_117 = data_d1[911:904];
        7'd115: vec_data_117 = data_d1[919:912];
        7'd116: vec_data_117 = data_d1[927:920];
        7'd117: vec_data_117 = data_d1[935:928];
        7'd118: vec_data_117 = data_d1[943:936];
    endcase
end

always @(
  vec_sum_118_d1
  or data_d1
  ) begin
    vec_data_118 = 8'b0;
    case(vec_sum_118_d1)
        7'd1: vec_data_118 = data_d1[7:0];
        7'd2: vec_data_118 = data_d1[15:8];
        7'd3: vec_data_118 = data_d1[23:16];
        7'd4: vec_data_118 = data_d1[31:24];
        7'd5: vec_data_118 = data_d1[39:32];
        7'd6: vec_data_118 = data_d1[47:40];
        7'd7: vec_data_118 = data_d1[55:48];
        7'd8: vec_data_118 = data_d1[63:56];
        7'd9: vec_data_118 = data_d1[71:64];
        7'd10: vec_data_118 = data_d1[79:72];
        7'd11: vec_data_118 = data_d1[87:80];
        7'd12: vec_data_118 = data_d1[95:88];
        7'd13: vec_data_118 = data_d1[103:96];
        7'd14: vec_data_118 = data_d1[111:104];
        7'd15: vec_data_118 = data_d1[119:112];
        7'd16: vec_data_118 = data_d1[127:120];
        7'd17: vec_data_118 = data_d1[135:128];
        7'd18: vec_data_118 = data_d1[143:136];
        7'd19: vec_data_118 = data_d1[151:144];
        7'd20: vec_data_118 = data_d1[159:152];
        7'd21: vec_data_118 = data_d1[167:160];
        7'd22: vec_data_118 = data_d1[175:168];
        7'd23: vec_data_118 = data_d1[183:176];
        7'd24: vec_data_118 = data_d1[191:184];
        7'd25: vec_data_118 = data_d1[199:192];
        7'd26: vec_data_118 = data_d1[207:200];
        7'd27: vec_data_118 = data_d1[215:208];
        7'd28: vec_data_118 = data_d1[223:216];
        7'd29: vec_data_118 = data_d1[231:224];
        7'd30: vec_data_118 = data_d1[239:232];
        7'd31: vec_data_118 = data_d1[247:240];
        7'd32: vec_data_118 = data_d1[255:248];
        7'd33: vec_data_118 = data_d1[263:256];
        7'd34: vec_data_118 = data_d1[271:264];
        7'd35: vec_data_118 = data_d1[279:272];
        7'd36: vec_data_118 = data_d1[287:280];
        7'd37: vec_data_118 = data_d1[295:288];
        7'd38: vec_data_118 = data_d1[303:296];
        7'd39: vec_data_118 = data_d1[311:304];
        7'd40: vec_data_118 = data_d1[319:312];
        7'd41: vec_data_118 = data_d1[327:320];
        7'd42: vec_data_118 = data_d1[335:328];
        7'd43: vec_data_118 = data_d1[343:336];
        7'd44: vec_data_118 = data_d1[351:344];
        7'd45: vec_data_118 = data_d1[359:352];
        7'd46: vec_data_118 = data_d1[367:360];
        7'd47: vec_data_118 = data_d1[375:368];
        7'd48: vec_data_118 = data_d1[383:376];
        7'd49: vec_data_118 = data_d1[391:384];
        7'd50: vec_data_118 = data_d1[399:392];
        7'd51: vec_data_118 = data_d1[407:400];
        7'd52: vec_data_118 = data_d1[415:408];
        7'd53: vec_data_118 = data_d1[423:416];
        7'd54: vec_data_118 = data_d1[431:424];
        7'd55: vec_data_118 = data_d1[439:432];
        7'd56: vec_data_118 = data_d1[447:440];
        7'd57: vec_data_118 = data_d1[455:448];
        7'd58: vec_data_118 = data_d1[463:456];
        7'd59: vec_data_118 = data_d1[471:464];
        7'd60: vec_data_118 = data_d1[479:472];
        7'd61: vec_data_118 = data_d1[487:480];
        7'd62: vec_data_118 = data_d1[495:488];
        7'd63: vec_data_118 = data_d1[503:496];
        7'd64: vec_data_118 = data_d1[511:504];
        7'd65: vec_data_118 = data_d1[519:512];
        7'd66: vec_data_118 = data_d1[527:520];
        7'd67: vec_data_118 = data_d1[535:528];
        7'd68: vec_data_118 = data_d1[543:536];
        7'd69: vec_data_118 = data_d1[551:544];
        7'd70: vec_data_118 = data_d1[559:552];
        7'd71: vec_data_118 = data_d1[567:560];
        7'd72: vec_data_118 = data_d1[575:568];
        7'd73: vec_data_118 = data_d1[583:576];
        7'd74: vec_data_118 = data_d1[591:584];
        7'd75: vec_data_118 = data_d1[599:592];
        7'd76: vec_data_118 = data_d1[607:600];
        7'd77: vec_data_118 = data_d1[615:608];
        7'd78: vec_data_118 = data_d1[623:616];
        7'd79: vec_data_118 = data_d1[631:624];
        7'd80: vec_data_118 = data_d1[639:632];
        7'd81: vec_data_118 = data_d1[647:640];
        7'd82: vec_data_118 = data_d1[655:648];
        7'd83: vec_data_118 = data_d1[663:656];
        7'd84: vec_data_118 = data_d1[671:664];
        7'd85: vec_data_118 = data_d1[679:672];
        7'd86: vec_data_118 = data_d1[687:680];
        7'd87: vec_data_118 = data_d1[695:688];
        7'd88: vec_data_118 = data_d1[703:696];
        7'd89: vec_data_118 = data_d1[711:704];
        7'd90: vec_data_118 = data_d1[719:712];
        7'd91: vec_data_118 = data_d1[727:720];
        7'd92: vec_data_118 = data_d1[735:728];
        7'd93: vec_data_118 = data_d1[743:736];
        7'd94: vec_data_118 = data_d1[751:744];
        7'd95: vec_data_118 = data_d1[759:752];
        7'd96: vec_data_118 = data_d1[767:760];
        7'd97: vec_data_118 = data_d1[775:768];
        7'd98: vec_data_118 = data_d1[783:776];
        7'd99: vec_data_118 = data_d1[791:784];
        7'd100: vec_data_118 = data_d1[799:792];
        7'd101: vec_data_118 = data_d1[807:800];
        7'd102: vec_data_118 = data_d1[815:808];
        7'd103: vec_data_118 = data_d1[823:816];
        7'd104: vec_data_118 = data_d1[831:824];
        7'd105: vec_data_118 = data_d1[839:832];
        7'd106: vec_data_118 = data_d1[847:840];
        7'd107: vec_data_118 = data_d1[855:848];
        7'd108: vec_data_118 = data_d1[863:856];
        7'd109: vec_data_118 = data_d1[871:864];
        7'd110: vec_data_118 = data_d1[879:872];
        7'd111: vec_data_118 = data_d1[887:880];
        7'd112: vec_data_118 = data_d1[895:888];
        7'd113: vec_data_118 = data_d1[903:896];
        7'd114: vec_data_118 = data_d1[911:904];
        7'd115: vec_data_118 = data_d1[919:912];
        7'd116: vec_data_118 = data_d1[927:920];
        7'd117: vec_data_118 = data_d1[935:928];
        7'd118: vec_data_118 = data_d1[943:936];
        7'd119: vec_data_118 = data_d1[951:944];
    endcase
end

always @(
  vec_sum_119_d1
  or data_d1
  ) begin
    vec_data_119 = 8'b0;
    case(vec_sum_119_d1)
        7'd1: vec_data_119 = data_d1[7:0];
        7'd2: vec_data_119 = data_d1[15:8];
        7'd3: vec_data_119 = data_d1[23:16];
        7'd4: vec_data_119 = data_d1[31:24];
        7'd5: vec_data_119 = data_d1[39:32];
        7'd6: vec_data_119 = data_d1[47:40];
        7'd7: vec_data_119 = data_d1[55:48];
        7'd8: vec_data_119 = data_d1[63:56];
        7'd9: vec_data_119 = data_d1[71:64];
        7'd10: vec_data_119 = data_d1[79:72];
        7'd11: vec_data_119 = data_d1[87:80];
        7'd12: vec_data_119 = data_d1[95:88];
        7'd13: vec_data_119 = data_d1[103:96];
        7'd14: vec_data_119 = data_d1[111:104];
        7'd15: vec_data_119 = data_d1[119:112];
        7'd16: vec_data_119 = data_d1[127:120];
        7'd17: vec_data_119 = data_d1[135:128];
        7'd18: vec_data_119 = data_d1[143:136];
        7'd19: vec_data_119 = data_d1[151:144];
        7'd20: vec_data_119 = data_d1[159:152];
        7'd21: vec_data_119 = data_d1[167:160];
        7'd22: vec_data_119 = data_d1[175:168];
        7'd23: vec_data_119 = data_d1[183:176];
        7'd24: vec_data_119 = data_d1[191:184];
        7'd25: vec_data_119 = data_d1[199:192];
        7'd26: vec_data_119 = data_d1[207:200];
        7'd27: vec_data_119 = data_d1[215:208];
        7'd28: vec_data_119 = data_d1[223:216];
        7'd29: vec_data_119 = data_d1[231:224];
        7'd30: vec_data_119 = data_d1[239:232];
        7'd31: vec_data_119 = data_d1[247:240];
        7'd32: vec_data_119 = data_d1[255:248];
        7'd33: vec_data_119 = data_d1[263:256];
        7'd34: vec_data_119 = data_d1[271:264];
        7'd35: vec_data_119 = data_d1[279:272];
        7'd36: vec_data_119 = data_d1[287:280];
        7'd37: vec_data_119 = data_d1[295:288];
        7'd38: vec_data_119 = data_d1[303:296];
        7'd39: vec_data_119 = data_d1[311:304];
        7'd40: vec_data_119 = data_d1[319:312];
        7'd41: vec_data_119 = data_d1[327:320];
        7'd42: vec_data_119 = data_d1[335:328];
        7'd43: vec_data_119 = data_d1[343:336];
        7'd44: vec_data_119 = data_d1[351:344];
        7'd45: vec_data_119 = data_d1[359:352];
        7'd46: vec_data_119 = data_d1[367:360];
        7'd47: vec_data_119 = data_d1[375:368];
        7'd48: vec_data_119 = data_d1[383:376];
        7'd49: vec_data_119 = data_d1[391:384];
        7'd50: vec_data_119 = data_d1[399:392];
        7'd51: vec_data_119 = data_d1[407:400];
        7'd52: vec_data_119 = data_d1[415:408];
        7'd53: vec_data_119 = data_d1[423:416];
        7'd54: vec_data_119 = data_d1[431:424];
        7'd55: vec_data_119 = data_d1[439:432];
        7'd56: vec_data_119 = data_d1[447:440];
        7'd57: vec_data_119 = data_d1[455:448];
        7'd58: vec_data_119 = data_d1[463:456];
        7'd59: vec_data_119 = data_d1[471:464];
        7'd60: vec_data_119 = data_d1[479:472];
        7'd61: vec_data_119 = data_d1[487:480];
        7'd62: vec_data_119 = data_d1[495:488];
        7'd63: vec_data_119 = data_d1[503:496];
        7'd64: vec_data_119 = data_d1[511:504];
        7'd65: vec_data_119 = data_d1[519:512];
        7'd66: vec_data_119 = data_d1[527:520];
        7'd67: vec_data_119 = data_d1[535:528];
        7'd68: vec_data_119 = data_d1[543:536];
        7'd69: vec_data_119 = data_d1[551:544];
        7'd70: vec_data_119 = data_d1[559:552];
        7'd71: vec_data_119 = data_d1[567:560];
        7'd72: vec_data_119 = data_d1[575:568];
        7'd73: vec_data_119 = data_d1[583:576];
        7'd74: vec_data_119 = data_d1[591:584];
        7'd75: vec_data_119 = data_d1[599:592];
        7'd76: vec_data_119 = data_d1[607:600];
        7'd77: vec_data_119 = data_d1[615:608];
        7'd78: vec_data_119 = data_d1[623:616];
        7'd79: vec_data_119 = data_d1[631:624];
        7'd80: vec_data_119 = data_d1[639:632];
        7'd81: vec_data_119 = data_d1[647:640];
        7'd82: vec_data_119 = data_d1[655:648];
        7'd83: vec_data_119 = data_d1[663:656];
        7'd84: vec_data_119 = data_d1[671:664];
        7'd85: vec_data_119 = data_d1[679:672];
        7'd86: vec_data_119 = data_d1[687:680];
        7'd87: vec_data_119 = data_d1[695:688];
        7'd88: vec_data_119 = data_d1[703:696];
        7'd89: vec_data_119 = data_d1[711:704];
        7'd90: vec_data_119 = data_d1[719:712];
        7'd91: vec_data_119 = data_d1[727:720];
        7'd92: vec_data_119 = data_d1[735:728];
        7'd93: vec_data_119 = data_d1[743:736];
        7'd94: vec_data_119 = data_d1[751:744];
        7'd95: vec_data_119 = data_d1[759:752];
        7'd96: vec_data_119 = data_d1[767:760];
        7'd97: vec_data_119 = data_d1[775:768];
        7'd98: vec_data_119 = data_d1[783:776];
        7'd99: vec_data_119 = data_d1[791:784];
        7'd100: vec_data_119 = data_d1[799:792];
        7'd101: vec_data_119 = data_d1[807:800];
        7'd102: vec_data_119 = data_d1[815:808];
        7'd103: vec_data_119 = data_d1[823:816];
        7'd104: vec_data_119 = data_d1[831:824];
        7'd105: vec_data_119 = data_d1[839:832];
        7'd106: vec_data_119 = data_d1[847:840];
        7'd107: vec_data_119 = data_d1[855:848];
        7'd108: vec_data_119 = data_d1[863:856];
        7'd109: vec_data_119 = data_d1[871:864];
        7'd110: vec_data_119 = data_d1[879:872];
        7'd111: vec_data_119 = data_d1[887:880];
        7'd112: vec_data_119 = data_d1[895:888];
        7'd113: vec_data_119 = data_d1[903:896];
        7'd114: vec_data_119 = data_d1[911:904];
        7'd115: vec_data_119 = data_d1[919:912];
        7'd116: vec_data_119 = data_d1[927:920];
        7'd117: vec_data_119 = data_d1[935:928];
        7'd118: vec_data_119 = data_d1[943:936];
        7'd119: vec_data_119 = data_d1[951:944];
        7'd120: vec_data_119 = data_d1[959:952];
    endcase
end

always @(
  vec_sum_120_d1
  or data_d1
  ) begin
    vec_data_120 = 8'b0;
    case(vec_sum_120_d1)
        7'd1: vec_data_120 = data_d1[7:0];
        7'd2: vec_data_120 = data_d1[15:8];
        7'd3: vec_data_120 = data_d1[23:16];
        7'd4: vec_data_120 = data_d1[31:24];
        7'd5: vec_data_120 = data_d1[39:32];
        7'd6: vec_data_120 = data_d1[47:40];
        7'd7: vec_data_120 = data_d1[55:48];
        7'd8: vec_data_120 = data_d1[63:56];
        7'd9: vec_data_120 = data_d1[71:64];
        7'd10: vec_data_120 = data_d1[79:72];
        7'd11: vec_data_120 = data_d1[87:80];
        7'd12: vec_data_120 = data_d1[95:88];
        7'd13: vec_data_120 = data_d1[103:96];
        7'd14: vec_data_120 = data_d1[111:104];
        7'd15: vec_data_120 = data_d1[119:112];
        7'd16: vec_data_120 = data_d1[127:120];
        7'd17: vec_data_120 = data_d1[135:128];
        7'd18: vec_data_120 = data_d1[143:136];
        7'd19: vec_data_120 = data_d1[151:144];
        7'd20: vec_data_120 = data_d1[159:152];
        7'd21: vec_data_120 = data_d1[167:160];
        7'd22: vec_data_120 = data_d1[175:168];
        7'd23: vec_data_120 = data_d1[183:176];
        7'd24: vec_data_120 = data_d1[191:184];
        7'd25: vec_data_120 = data_d1[199:192];
        7'd26: vec_data_120 = data_d1[207:200];
        7'd27: vec_data_120 = data_d1[215:208];
        7'd28: vec_data_120 = data_d1[223:216];
        7'd29: vec_data_120 = data_d1[231:224];
        7'd30: vec_data_120 = data_d1[239:232];
        7'd31: vec_data_120 = data_d1[247:240];
        7'd32: vec_data_120 = data_d1[255:248];
        7'd33: vec_data_120 = data_d1[263:256];
        7'd34: vec_data_120 = data_d1[271:264];
        7'd35: vec_data_120 = data_d1[279:272];
        7'd36: vec_data_120 = data_d1[287:280];
        7'd37: vec_data_120 = data_d1[295:288];
        7'd38: vec_data_120 = data_d1[303:296];
        7'd39: vec_data_120 = data_d1[311:304];
        7'd40: vec_data_120 = data_d1[319:312];
        7'd41: vec_data_120 = data_d1[327:320];
        7'd42: vec_data_120 = data_d1[335:328];
        7'd43: vec_data_120 = data_d1[343:336];
        7'd44: vec_data_120 = data_d1[351:344];
        7'd45: vec_data_120 = data_d1[359:352];
        7'd46: vec_data_120 = data_d1[367:360];
        7'd47: vec_data_120 = data_d1[375:368];
        7'd48: vec_data_120 = data_d1[383:376];
        7'd49: vec_data_120 = data_d1[391:384];
        7'd50: vec_data_120 = data_d1[399:392];
        7'd51: vec_data_120 = data_d1[407:400];
        7'd52: vec_data_120 = data_d1[415:408];
        7'd53: vec_data_120 = data_d1[423:416];
        7'd54: vec_data_120 = data_d1[431:424];
        7'd55: vec_data_120 = data_d1[439:432];
        7'd56: vec_data_120 = data_d1[447:440];
        7'd57: vec_data_120 = data_d1[455:448];
        7'd58: vec_data_120 = data_d1[463:456];
        7'd59: vec_data_120 = data_d1[471:464];
        7'd60: vec_data_120 = data_d1[479:472];
        7'd61: vec_data_120 = data_d1[487:480];
        7'd62: vec_data_120 = data_d1[495:488];
        7'd63: vec_data_120 = data_d1[503:496];
        7'd64: vec_data_120 = data_d1[511:504];
        7'd65: vec_data_120 = data_d1[519:512];
        7'd66: vec_data_120 = data_d1[527:520];
        7'd67: vec_data_120 = data_d1[535:528];
        7'd68: vec_data_120 = data_d1[543:536];
        7'd69: vec_data_120 = data_d1[551:544];
        7'd70: vec_data_120 = data_d1[559:552];
        7'd71: vec_data_120 = data_d1[567:560];
        7'd72: vec_data_120 = data_d1[575:568];
        7'd73: vec_data_120 = data_d1[583:576];
        7'd74: vec_data_120 = data_d1[591:584];
        7'd75: vec_data_120 = data_d1[599:592];
        7'd76: vec_data_120 = data_d1[607:600];
        7'd77: vec_data_120 = data_d1[615:608];
        7'd78: vec_data_120 = data_d1[623:616];
        7'd79: vec_data_120 = data_d1[631:624];
        7'd80: vec_data_120 = data_d1[639:632];
        7'd81: vec_data_120 = data_d1[647:640];
        7'd82: vec_data_120 = data_d1[655:648];
        7'd83: vec_data_120 = data_d1[663:656];
        7'd84: vec_data_120 = data_d1[671:664];
        7'd85: vec_data_120 = data_d1[679:672];
        7'd86: vec_data_120 = data_d1[687:680];
        7'd87: vec_data_120 = data_d1[695:688];
        7'd88: vec_data_120 = data_d1[703:696];
        7'd89: vec_data_120 = data_d1[711:704];
        7'd90: vec_data_120 = data_d1[719:712];
        7'd91: vec_data_120 = data_d1[727:720];
        7'd92: vec_data_120 = data_d1[735:728];
        7'd93: vec_data_120 = data_d1[743:736];
        7'd94: vec_data_120 = data_d1[751:744];
        7'd95: vec_data_120 = data_d1[759:752];
        7'd96: vec_data_120 = data_d1[767:760];
        7'd97: vec_data_120 = data_d1[775:768];
        7'd98: vec_data_120 = data_d1[783:776];
        7'd99: vec_data_120 = data_d1[791:784];
        7'd100: vec_data_120 = data_d1[799:792];
        7'd101: vec_data_120 = data_d1[807:800];
        7'd102: vec_data_120 = data_d1[815:808];
        7'd103: vec_data_120 = data_d1[823:816];
        7'd104: vec_data_120 = data_d1[831:824];
        7'd105: vec_data_120 = data_d1[839:832];
        7'd106: vec_data_120 = data_d1[847:840];
        7'd107: vec_data_120 = data_d1[855:848];
        7'd108: vec_data_120 = data_d1[863:856];
        7'd109: vec_data_120 = data_d1[871:864];
        7'd110: vec_data_120 = data_d1[879:872];
        7'd111: vec_data_120 = data_d1[887:880];
        7'd112: vec_data_120 = data_d1[895:888];
        7'd113: vec_data_120 = data_d1[903:896];
        7'd114: vec_data_120 = data_d1[911:904];
        7'd115: vec_data_120 = data_d1[919:912];
        7'd116: vec_data_120 = data_d1[927:920];
        7'd117: vec_data_120 = data_d1[935:928];
        7'd118: vec_data_120 = data_d1[943:936];
        7'd119: vec_data_120 = data_d1[951:944];
        7'd120: vec_data_120 = data_d1[959:952];
        7'd121: vec_data_120 = data_d1[967:960];
    endcase
end

always @(
  vec_sum_121_d1
  or data_d1
  ) begin
    vec_data_121 = 8'b0;
    case(vec_sum_121_d1)
        7'd1: vec_data_121 = data_d1[7:0];
        7'd2: vec_data_121 = data_d1[15:8];
        7'd3: vec_data_121 = data_d1[23:16];
        7'd4: vec_data_121 = data_d1[31:24];
        7'd5: vec_data_121 = data_d1[39:32];
        7'd6: vec_data_121 = data_d1[47:40];
        7'd7: vec_data_121 = data_d1[55:48];
        7'd8: vec_data_121 = data_d1[63:56];
        7'd9: vec_data_121 = data_d1[71:64];
        7'd10: vec_data_121 = data_d1[79:72];
        7'd11: vec_data_121 = data_d1[87:80];
        7'd12: vec_data_121 = data_d1[95:88];
        7'd13: vec_data_121 = data_d1[103:96];
        7'd14: vec_data_121 = data_d1[111:104];
        7'd15: vec_data_121 = data_d1[119:112];
        7'd16: vec_data_121 = data_d1[127:120];
        7'd17: vec_data_121 = data_d1[135:128];
        7'd18: vec_data_121 = data_d1[143:136];
        7'd19: vec_data_121 = data_d1[151:144];
        7'd20: vec_data_121 = data_d1[159:152];
        7'd21: vec_data_121 = data_d1[167:160];
        7'd22: vec_data_121 = data_d1[175:168];
        7'd23: vec_data_121 = data_d1[183:176];
        7'd24: vec_data_121 = data_d1[191:184];
        7'd25: vec_data_121 = data_d1[199:192];
        7'd26: vec_data_121 = data_d1[207:200];
        7'd27: vec_data_121 = data_d1[215:208];
        7'd28: vec_data_121 = data_d1[223:216];
        7'd29: vec_data_121 = data_d1[231:224];
        7'd30: vec_data_121 = data_d1[239:232];
        7'd31: vec_data_121 = data_d1[247:240];
        7'd32: vec_data_121 = data_d1[255:248];
        7'd33: vec_data_121 = data_d1[263:256];
        7'd34: vec_data_121 = data_d1[271:264];
        7'd35: vec_data_121 = data_d1[279:272];
        7'd36: vec_data_121 = data_d1[287:280];
        7'd37: vec_data_121 = data_d1[295:288];
        7'd38: vec_data_121 = data_d1[303:296];
        7'd39: vec_data_121 = data_d1[311:304];
        7'd40: vec_data_121 = data_d1[319:312];
        7'd41: vec_data_121 = data_d1[327:320];
        7'd42: vec_data_121 = data_d1[335:328];
        7'd43: vec_data_121 = data_d1[343:336];
        7'd44: vec_data_121 = data_d1[351:344];
        7'd45: vec_data_121 = data_d1[359:352];
        7'd46: vec_data_121 = data_d1[367:360];
        7'd47: vec_data_121 = data_d1[375:368];
        7'd48: vec_data_121 = data_d1[383:376];
        7'd49: vec_data_121 = data_d1[391:384];
        7'd50: vec_data_121 = data_d1[399:392];
        7'd51: vec_data_121 = data_d1[407:400];
        7'd52: vec_data_121 = data_d1[415:408];
        7'd53: vec_data_121 = data_d1[423:416];
        7'd54: vec_data_121 = data_d1[431:424];
        7'd55: vec_data_121 = data_d1[439:432];
        7'd56: vec_data_121 = data_d1[447:440];
        7'd57: vec_data_121 = data_d1[455:448];
        7'd58: vec_data_121 = data_d1[463:456];
        7'd59: vec_data_121 = data_d1[471:464];
        7'd60: vec_data_121 = data_d1[479:472];
        7'd61: vec_data_121 = data_d1[487:480];
        7'd62: vec_data_121 = data_d1[495:488];
        7'd63: vec_data_121 = data_d1[503:496];
        7'd64: vec_data_121 = data_d1[511:504];
        7'd65: vec_data_121 = data_d1[519:512];
        7'd66: vec_data_121 = data_d1[527:520];
        7'd67: vec_data_121 = data_d1[535:528];
        7'd68: vec_data_121 = data_d1[543:536];
        7'd69: vec_data_121 = data_d1[551:544];
        7'd70: vec_data_121 = data_d1[559:552];
        7'd71: vec_data_121 = data_d1[567:560];
        7'd72: vec_data_121 = data_d1[575:568];
        7'd73: vec_data_121 = data_d1[583:576];
        7'd74: vec_data_121 = data_d1[591:584];
        7'd75: vec_data_121 = data_d1[599:592];
        7'd76: vec_data_121 = data_d1[607:600];
        7'd77: vec_data_121 = data_d1[615:608];
        7'd78: vec_data_121 = data_d1[623:616];
        7'd79: vec_data_121 = data_d1[631:624];
        7'd80: vec_data_121 = data_d1[639:632];
        7'd81: vec_data_121 = data_d1[647:640];
        7'd82: vec_data_121 = data_d1[655:648];
        7'd83: vec_data_121 = data_d1[663:656];
        7'd84: vec_data_121 = data_d1[671:664];
        7'd85: vec_data_121 = data_d1[679:672];
        7'd86: vec_data_121 = data_d1[687:680];
        7'd87: vec_data_121 = data_d1[695:688];
        7'd88: vec_data_121 = data_d1[703:696];
        7'd89: vec_data_121 = data_d1[711:704];
        7'd90: vec_data_121 = data_d1[719:712];
        7'd91: vec_data_121 = data_d1[727:720];
        7'd92: vec_data_121 = data_d1[735:728];
        7'd93: vec_data_121 = data_d1[743:736];
        7'd94: vec_data_121 = data_d1[751:744];
        7'd95: vec_data_121 = data_d1[759:752];
        7'd96: vec_data_121 = data_d1[767:760];
        7'd97: vec_data_121 = data_d1[775:768];
        7'd98: vec_data_121 = data_d1[783:776];
        7'd99: vec_data_121 = data_d1[791:784];
        7'd100: vec_data_121 = data_d1[799:792];
        7'd101: vec_data_121 = data_d1[807:800];
        7'd102: vec_data_121 = data_d1[815:808];
        7'd103: vec_data_121 = data_d1[823:816];
        7'd104: vec_data_121 = data_d1[831:824];
        7'd105: vec_data_121 = data_d1[839:832];
        7'd106: vec_data_121 = data_d1[847:840];
        7'd107: vec_data_121 = data_d1[855:848];
        7'd108: vec_data_121 = data_d1[863:856];
        7'd109: vec_data_121 = data_d1[871:864];
        7'd110: vec_data_121 = data_d1[879:872];
        7'd111: vec_data_121 = data_d1[887:880];
        7'd112: vec_data_121 = data_d1[895:888];
        7'd113: vec_data_121 = data_d1[903:896];
        7'd114: vec_data_121 = data_d1[911:904];
        7'd115: vec_data_121 = data_d1[919:912];
        7'd116: vec_data_121 = data_d1[927:920];
        7'd117: vec_data_121 = data_d1[935:928];
        7'd118: vec_data_121 = data_d1[943:936];
        7'd119: vec_data_121 = data_d1[951:944];
        7'd120: vec_data_121 = data_d1[959:952];
        7'd121: vec_data_121 = data_d1[967:960];
        7'd122: vec_data_121 = data_d1[975:968];
    endcase
end

always @(
  vec_sum_122_d1
  or data_d1
  ) begin
    vec_data_122 = 8'b0;
    case(vec_sum_122_d1)
        7'd1: vec_data_122 = data_d1[7:0];
        7'd2: vec_data_122 = data_d1[15:8];
        7'd3: vec_data_122 = data_d1[23:16];
        7'd4: vec_data_122 = data_d1[31:24];
        7'd5: vec_data_122 = data_d1[39:32];
        7'd6: vec_data_122 = data_d1[47:40];
        7'd7: vec_data_122 = data_d1[55:48];
        7'd8: vec_data_122 = data_d1[63:56];
        7'd9: vec_data_122 = data_d1[71:64];
        7'd10: vec_data_122 = data_d1[79:72];
        7'd11: vec_data_122 = data_d1[87:80];
        7'd12: vec_data_122 = data_d1[95:88];
        7'd13: vec_data_122 = data_d1[103:96];
        7'd14: vec_data_122 = data_d1[111:104];
        7'd15: vec_data_122 = data_d1[119:112];
        7'd16: vec_data_122 = data_d1[127:120];
        7'd17: vec_data_122 = data_d1[135:128];
        7'd18: vec_data_122 = data_d1[143:136];
        7'd19: vec_data_122 = data_d1[151:144];
        7'd20: vec_data_122 = data_d1[159:152];
        7'd21: vec_data_122 = data_d1[167:160];
        7'd22: vec_data_122 = data_d1[175:168];
        7'd23: vec_data_122 = data_d1[183:176];
        7'd24: vec_data_122 = data_d1[191:184];
        7'd25: vec_data_122 = data_d1[199:192];
        7'd26: vec_data_122 = data_d1[207:200];
        7'd27: vec_data_122 = data_d1[215:208];
        7'd28: vec_data_122 = data_d1[223:216];
        7'd29: vec_data_122 = data_d1[231:224];
        7'd30: vec_data_122 = data_d1[239:232];
        7'd31: vec_data_122 = data_d1[247:240];
        7'd32: vec_data_122 = data_d1[255:248];
        7'd33: vec_data_122 = data_d1[263:256];
        7'd34: vec_data_122 = data_d1[271:264];
        7'd35: vec_data_122 = data_d1[279:272];
        7'd36: vec_data_122 = data_d1[287:280];
        7'd37: vec_data_122 = data_d1[295:288];
        7'd38: vec_data_122 = data_d1[303:296];
        7'd39: vec_data_122 = data_d1[311:304];
        7'd40: vec_data_122 = data_d1[319:312];
        7'd41: vec_data_122 = data_d1[327:320];
        7'd42: vec_data_122 = data_d1[335:328];
        7'd43: vec_data_122 = data_d1[343:336];
        7'd44: vec_data_122 = data_d1[351:344];
        7'd45: vec_data_122 = data_d1[359:352];
        7'd46: vec_data_122 = data_d1[367:360];
        7'd47: vec_data_122 = data_d1[375:368];
        7'd48: vec_data_122 = data_d1[383:376];
        7'd49: vec_data_122 = data_d1[391:384];
        7'd50: vec_data_122 = data_d1[399:392];
        7'd51: vec_data_122 = data_d1[407:400];
        7'd52: vec_data_122 = data_d1[415:408];
        7'd53: vec_data_122 = data_d1[423:416];
        7'd54: vec_data_122 = data_d1[431:424];
        7'd55: vec_data_122 = data_d1[439:432];
        7'd56: vec_data_122 = data_d1[447:440];
        7'd57: vec_data_122 = data_d1[455:448];
        7'd58: vec_data_122 = data_d1[463:456];
        7'd59: vec_data_122 = data_d1[471:464];
        7'd60: vec_data_122 = data_d1[479:472];
        7'd61: vec_data_122 = data_d1[487:480];
        7'd62: vec_data_122 = data_d1[495:488];
        7'd63: vec_data_122 = data_d1[503:496];
        7'd64: vec_data_122 = data_d1[511:504];
        7'd65: vec_data_122 = data_d1[519:512];
        7'd66: vec_data_122 = data_d1[527:520];
        7'd67: vec_data_122 = data_d1[535:528];
        7'd68: vec_data_122 = data_d1[543:536];
        7'd69: vec_data_122 = data_d1[551:544];
        7'd70: vec_data_122 = data_d1[559:552];
        7'd71: vec_data_122 = data_d1[567:560];
        7'd72: vec_data_122 = data_d1[575:568];
        7'd73: vec_data_122 = data_d1[583:576];
        7'd74: vec_data_122 = data_d1[591:584];
        7'd75: vec_data_122 = data_d1[599:592];
        7'd76: vec_data_122 = data_d1[607:600];
        7'd77: vec_data_122 = data_d1[615:608];
        7'd78: vec_data_122 = data_d1[623:616];
        7'd79: vec_data_122 = data_d1[631:624];
        7'd80: vec_data_122 = data_d1[639:632];
        7'd81: vec_data_122 = data_d1[647:640];
        7'd82: vec_data_122 = data_d1[655:648];
        7'd83: vec_data_122 = data_d1[663:656];
        7'd84: vec_data_122 = data_d1[671:664];
        7'd85: vec_data_122 = data_d1[679:672];
        7'd86: vec_data_122 = data_d1[687:680];
        7'd87: vec_data_122 = data_d1[695:688];
        7'd88: vec_data_122 = data_d1[703:696];
        7'd89: vec_data_122 = data_d1[711:704];
        7'd90: vec_data_122 = data_d1[719:712];
        7'd91: vec_data_122 = data_d1[727:720];
        7'd92: vec_data_122 = data_d1[735:728];
        7'd93: vec_data_122 = data_d1[743:736];
        7'd94: vec_data_122 = data_d1[751:744];
        7'd95: vec_data_122 = data_d1[759:752];
        7'd96: vec_data_122 = data_d1[767:760];
        7'd97: vec_data_122 = data_d1[775:768];
        7'd98: vec_data_122 = data_d1[783:776];
        7'd99: vec_data_122 = data_d1[791:784];
        7'd100: vec_data_122 = data_d1[799:792];
        7'd101: vec_data_122 = data_d1[807:800];
        7'd102: vec_data_122 = data_d1[815:808];
        7'd103: vec_data_122 = data_d1[823:816];
        7'd104: vec_data_122 = data_d1[831:824];
        7'd105: vec_data_122 = data_d1[839:832];
        7'd106: vec_data_122 = data_d1[847:840];
        7'd107: vec_data_122 = data_d1[855:848];
        7'd108: vec_data_122 = data_d1[863:856];
        7'd109: vec_data_122 = data_d1[871:864];
        7'd110: vec_data_122 = data_d1[879:872];
        7'd111: vec_data_122 = data_d1[887:880];
        7'd112: vec_data_122 = data_d1[895:888];
        7'd113: vec_data_122 = data_d1[903:896];
        7'd114: vec_data_122 = data_d1[911:904];
        7'd115: vec_data_122 = data_d1[919:912];
        7'd116: vec_data_122 = data_d1[927:920];
        7'd117: vec_data_122 = data_d1[935:928];
        7'd118: vec_data_122 = data_d1[943:936];
        7'd119: vec_data_122 = data_d1[951:944];
        7'd120: vec_data_122 = data_d1[959:952];
        7'd121: vec_data_122 = data_d1[967:960];
        7'd122: vec_data_122 = data_d1[975:968];
        7'd123: vec_data_122 = data_d1[983:976];
    endcase
end

always @(
  vec_sum_123_d1
  or data_d1
  ) begin
    vec_data_123 = 8'b0;
    case(vec_sum_123_d1)
        7'd1: vec_data_123 = data_d1[7:0];
        7'd2: vec_data_123 = data_d1[15:8];
        7'd3: vec_data_123 = data_d1[23:16];
        7'd4: vec_data_123 = data_d1[31:24];
        7'd5: vec_data_123 = data_d1[39:32];
        7'd6: vec_data_123 = data_d1[47:40];
        7'd7: vec_data_123 = data_d1[55:48];
        7'd8: vec_data_123 = data_d1[63:56];
        7'd9: vec_data_123 = data_d1[71:64];
        7'd10: vec_data_123 = data_d1[79:72];
        7'd11: vec_data_123 = data_d1[87:80];
        7'd12: vec_data_123 = data_d1[95:88];
        7'd13: vec_data_123 = data_d1[103:96];
        7'd14: vec_data_123 = data_d1[111:104];
        7'd15: vec_data_123 = data_d1[119:112];
        7'd16: vec_data_123 = data_d1[127:120];
        7'd17: vec_data_123 = data_d1[135:128];
        7'd18: vec_data_123 = data_d1[143:136];
        7'd19: vec_data_123 = data_d1[151:144];
        7'd20: vec_data_123 = data_d1[159:152];
        7'd21: vec_data_123 = data_d1[167:160];
        7'd22: vec_data_123 = data_d1[175:168];
        7'd23: vec_data_123 = data_d1[183:176];
        7'd24: vec_data_123 = data_d1[191:184];
        7'd25: vec_data_123 = data_d1[199:192];
        7'd26: vec_data_123 = data_d1[207:200];
        7'd27: vec_data_123 = data_d1[215:208];
        7'd28: vec_data_123 = data_d1[223:216];
        7'd29: vec_data_123 = data_d1[231:224];
        7'd30: vec_data_123 = data_d1[239:232];
        7'd31: vec_data_123 = data_d1[247:240];
        7'd32: vec_data_123 = data_d1[255:248];
        7'd33: vec_data_123 = data_d1[263:256];
        7'd34: vec_data_123 = data_d1[271:264];
        7'd35: vec_data_123 = data_d1[279:272];
        7'd36: vec_data_123 = data_d1[287:280];
        7'd37: vec_data_123 = data_d1[295:288];
        7'd38: vec_data_123 = data_d1[303:296];
        7'd39: vec_data_123 = data_d1[311:304];
        7'd40: vec_data_123 = data_d1[319:312];
        7'd41: vec_data_123 = data_d1[327:320];
        7'd42: vec_data_123 = data_d1[335:328];
        7'd43: vec_data_123 = data_d1[343:336];
        7'd44: vec_data_123 = data_d1[351:344];
        7'd45: vec_data_123 = data_d1[359:352];
        7'd46: vec_data_123 = data_d1[367:360];
        7'd47: vec_data_123 = data_d1[375:368];
        7'd48: vec_data_123 = data_d1[383:376];
        7'd49: vec_data_123 = data_d1[391:384];
        7'd50: vec_data_123 = data_d1[399:392];
        7'd51: vec_data_123 = data_d1[407:400];
        7'd52: vec_data_123 = data_d1[415:408];
        7'd53: vec_data_123 = data_d1[423:416];
        7'd54: vec_data_123 = data_d1[431:424];
        7'd55: vec_data_123 = data_d1[439:432];
        7'd56: vec_data_123 = data_d1[447:440];
        7'd57: vec_data_123 = data_d1[455:448];
        7'd58: vec_data_123 = data_d1[463:456];
        7'd59: vec_data_123 = data_d1[471:464];
        7'd60: vec_data_123 = data_d1[479:472];
        7'd61: vec_data_123 = data_d1[487:480];
        7'd62: vec_data_123 = data_d1[495:488];
        7'd63: vec_data_123 = data_d1[503:496];
        7'd64: vec_data_123 = data_d1[511:504];
        7'd65: vec_data_123 = data_d1[519:512];
        7'd66: vec_data_123 = data_d1[527:520];
        7'd67: vec_data_123 = data_d1[535:528];
        7'd68: vec_data_123 = data_d1[543:536];
        7'd69: vec_data_123 = data_d1[551:544];
        7'd70: vec_data_123 = data_d1[559:552];
        7'd71: vec_data_123 = data_d1[567:560];
        7'd72: vec_data_123 = data_d1[575:568];
        7'd73: vec_data_123 = data_d1[583:576];
        7'd74: vec_data_123 = data_d1[591:584];
        7'd75: vec_data_123 = data_d1[599:592];
        7'd76: vec_data_123 = data_d1[607:600];
        7'd77: vec_data_123 = data_d1[615:608];
        7'd78: vec_data_123 = data_d1[623:616];
        7'd79: vec_data_123 = data_d1[631:624];
        7'd80: vec_data_123 = data_d1[639:632];
        7'd81: vec_data_123 = data_d1[647:640];
        7'd82: vec_data_123 = data_d1[655:648];
        7'd83: vec_data_123 = data_d1[663:656];
        7'd84: vec_data_123 = data_d1[671:664];
        7'd85: vec_data_123 = data_d1[679:672];
        7'd86: vec_data_123 = data_d1[687:680];
        7'd87: vec_data_123 = data_d1[695:688];
        7'd88: vec_data_123 = data_d1[703:696];
        7'd89: vec_data_123 = data_d1[711:704];
        7'd90: vec_data_123 = data_d1[719:712];
        7'd91: vec_data_123 = data_d1[727:720];
        7'd92: vec_data_123 = data_d1[735:728];
        7'd93: vec_data_123 = data_d1[743:736];
        7'd94: vec_data_123 = data_d1[751:744];
        7'd95: vec_data_123 = data_d1[759:752];
        7'd96: vec_data_123 = data_d1[767:760];
        7'd97: vec_data_123 = data_d1[775:768];
        7'd98: vec_data_123 = data_d1[783:776];
        7'd99: vec_data_123 = data_d1[791:784];
        7'd100: vec_data_123 = data_d1[799:792];
        7'd101: vec_data_123 = data_d1[807:800];
        7'd102: vec_data_123 = data_d1[815:808];
        7'd103: vec_data_123 = data_d1[823:816];
        7'd104: vec_data_123 = data_d1[831:824];
        7'd105: vec_data_123 = data_d1[839:832];
        7'd106: vec_data_123 = data_d1[847:840];
        7'd107: vec_data_123 = data_d1[855:848];
        7'd108: vec_data_123 = data_d1[863:856];
        7'd109: vec_data_123 = data_d1[871:864];
        7'd110: vec_data_123 = data_d1[879:872];
        7'd111: vec_data_123 = data_d1[887:880];
        7'd112: vec_data_123 = data_d1[895:888];
        7'd113: vec_data_123 = data_d1[903:896];
        7'd114: vec_data_123 = data_d1[911:904];
        7'd115: vec_data_123 = data_d1[919:912];
        7'd116: vec_data_123 = data_d1[927:920];
        7'd117: vec_data_123 = data_d1[935:928];
        7'd118: vec_data_123 = data_d1[943:936];
        7'd119: vec_data_123 = data_d1[951:944];
        7'd120: vec_data_123 = data_d1[959:952];
        7'd121: vec_data_123 = data_d1[967:960];
        7'd122: vec_data_123 = data_d1[975:968];
        7'd123: vec_data_123 = data_d1[983:976];
        7'd124: vec_data_123 = data_d1[991:984];
    endcase
end

always @(
  vec_sum_124_d1
  or data_d1
  ) begin
    vec_data_124 = 8'b0;
    case(vec_sum_124_d1)
        7'd1: vec_data_124 = data_d1[7:0];
        7'd2: vec_data_124 = data_d1[15:8];
        7'd3: vec_data_124 = data_d1[23:16];
        7'd4: vec_data_124 = data_d1[31:24];
        7'd5: vec_data_124 = data_d1[39:32];
        7'd6: vec_data_124 = data_d1[47:40];
        7'd7: vec_data_124 = data_d1[55:48];
        7'd8: vec_data_124 = data_d1[63:56];
        7'd9: vec_data_124 = data_d1[71:64];
        7'd10: vec_data_124 = data_d1[79:72];
        7'd11: vec_data_124 = data_d1[87:80];
        7'd12: vec_data_124 = data_d1[95:88];
        7'd13: vec_data_124 = data_d1[103:96];
        7'd14: vec_data_124 = data_d1[111:104];
        7'd15: vec_data_124 = data_d1[119:112];
        7'd16: vec_data_124 = data_d1[127:120];
        7'd17: vec_data_124 = data_d1[135:128];
        7'd18: vec_data_124 = data_d1[143:136];
        7'd19: vec_data_124 = data_d1[151:144];
        7'd20: vec_data_124 = data_d1[159:152];
        7'd21: vec_data_124 = data_d1[167:160];
        7'd22: vec_data_124 = data_d1[175:168];
        7'd23: vec_data_124 = data_d1[183:176];
        7'd24: vec_data_124 = data_d1[191:184];
        7'd25: vec_data_124 = data_d1[199:192];
        7'd26: vec_data_124 = data_d1[207:200];
        7'd27: vec_data_124 = data_d1[215:208];
        7'd28: vec_data_124 = data_d1[223:216];
        7'd29: vec_data_124 = data_d1[231:224];
        7'd30: vec_data_124 = data_d1[239:232];
        7'd31: vec_data_124 = data_d1[247:240];
        7'd32: vec_data_124 = data_d1[255:248];
        7'd33: vec_data_124 = data_d1[263:256];
        7'd34: vec_data_124 = data_d1[271:264];
        7'd35: vec_data_124 = data_d1[279:272];
        7'd36: vec_data_124 = data_d1[287:280];
        7'd37: vec_data_124 = data_d1[295:288];
        7'd38: vec_data_124 = data_d1[303:296];
        7'd39: vec_data_124 = data_d1[311:304];
        7'd40: vec_data_124 = data_d1[319:312];
        7'd41: vec_data_124 = data_d1[327:320];
        7'd42: vec_data_124 = data_d1[335:328];
        7'd43: vec_data_124 = data_d1[343:336];
        7'd44: vec_data_124 = data_d1[351:344];
        7'd45: vec_data_124 = data_d1[359:352];
        7'd46: vec_data_124 = data_d1[367:360];
        7'd47: vec_data_124 = data_d1[375:368];
        7'd48: vec_data_124 = data_d1[383:376];
        7'd49: vec_data_124 = data_d1[391:384];
        7'd50: vec_data_124 = data_d1[399:392];
        7'd51: vec_data_124 = data_d1[407:400];
        7'd52: vec_data_124 = data_d1[415:408];
        7'd53: vec_data_124 = data_d1[423:416];
        7'd54: vec_data_124 = data_d1[431:424];
        7'd55: vec_data_124 = data_d1[439:432];
        7'd56: vec_data_124 = data_d1[447:440];
        7'd57: vec_data_124 = data_d1[455:448];
        7'd58: vec_data_124 = data_d1[463:456];
        7'd59: vec_data_124 = data_d1[471:464];
        7'd60: vec_data_124 = data_d1[479:472];
        7'd61: vec_data_124 = data_d1[487:480];
        7'd62: vec_data_124 = data_d1[495:488];
        7'd63: vec_data_124 = data_d1[503:496];
        7'd64: vec_data_124 = data_d1[511:504];
        7'd65: vec_data_124 = data_d1[519:512];
        7'd66: vec_data_124 = data_d1[527:520];
        7'd67: vec_data_124 = data_d1[535:528];
        7'd68: vec_data_124 = data_d1[543:536];
        7'd69: vec_data_124 = data_d1[551:544];
        7'd70: vec_data_124 = data_d1[559:552];
        7'd71: vec_data_124 = data_d1[567:560];
        7'd72: vec_data_124 = data_d1[575:568];
        7'd73: vec_data_124 = data_d1[583:576];
        7'd74: vec_data_124 = data_d1[591:584];
        7'd75: vec_data_124 = data_d1[599:592];
        7'd76: vec_data_124 = data_d1[607:600];
        7'd77: vec_data_124 = data_d1[615:608];
        7'd78: vec_data_124 = data_d1[623:616];
        7'd79: vec_data_124 = data_d1[631:624];
        7'd80: vec_data_124 = data_d1[639:632];
        7'd81: vec_data_124 = data_d1[647:640];
        7'd82: vec_data_124 = data_d1[655:648];
        7'd83: vec_data_124 = data_d1[663:656];
        7'd84: vec_data_124 = data_d1[671:664];
        7'd85: vec_data_124 = data_d1[679:672];
        7'd86: vec_data_124 = data_d1[687:680];
        7'd87: vec_data_124 = data_d1[695:688];
        7'd88: vec_data_124 = data_d1[703:696];
        7'd89: vec_data_124 = data_d1[711:704];
        7'd90: vec_data_124 = data_d1[719:712];
        7'd91: vec_data_124 = data_d1[727:720];
        7'd92: vec_data_124 = data_d1[735:728];
        7'd93: vec_data_124 = data_d1[743:736];
        7'd94: vec_data_124 = data_d1[751:744];
        7'd95: vec_data_124 = data_d1[759:752];
        7'd96: vec_data_124 = data_d1[767:760];
        7'd97: vec_data_124 = data_d1[775:768];
        7'd98: vec_data_124 = data_d1[783:776];
        7'd99: vec_data_124 = data_d1[791:784];
        7'd100: vec_data_124 = data_d1[799:792];
        7'd101: vec_data_124 = data_d1[807:800];
        7'd102: vec_data_124 = data_d1[815:808];
        7'd103: vec_data_124 = data_d1[823:816];
        7'd104: vec_data_124 = data_d1[831:824];
        7'd105: vec_data_124 = data_d1[839:832];
        7'd106: vec_data_124 = data_d1[847:840];
        7'd107: vec_data_124 = data_d1[855:848];
        7'd108: vec_data_124 = data_d1[863:856];
        7'd109: vec_data_124 = data_d1[871:864];
        7'd110: vec_data_124 = data_d1[879:872];
        7'd111: vec_data_124 = data_d1[887:880];
        7'd112: vec_data_124 = data_d1[895:888];
        7'd113: vec_data_124 = data_d1[903:896];
        7'd114: vec_data_124 = data_d1[911:904];
        7'd115: vec_data_124 = data_d1[919:912];
        7'd116: vec_data_124 = data_d1[927:920];
        7'd117: vec_data_124 = data_d1[935:928];
        7'd118: vec_data_124 = data_d1[943:936];
        7'd119: vec_data_124 = data_d1[951:944];
        7'd120: vec_data_124 = data_d1[959:952];
        7'd121: vec_data_124 = data_d1[967:960];
        7'd122: vec_data_124 = data_d1[975:968];
        7'd123: vec_data_124 = data_d1[983:976];
        7'd124: vec_data_124 = data_d1[991:984];
        7'd125: vec_data_124 = data_d1[999:992];
    endcase
end

always @(
  vec_sum_125_d1
  or data_d1
  ) begin
    vec_data_125 = 8'b0;
    case(vec_sum_125_d1)
        7'd1: vec_data_125 = data_d1[7:0];
        7'd2: vec_data_125 = data_d1[15:8];
        7'd3: vec_data_125 = data_d1[23:16];
        7'd4: vec_data_125 = data_d1[31:24];
        7'd5: vec_data_125 = data_d1[39:32];
        7'd6: vec_data_125 = data_d1[47:40];
        7'd7: vec_data_125 = data_d1[55:48];
        7'd8: vec_data_125 = data_d1[63:56];
        7'd9: vec_data_125 = data_d1[71:64];
        7'd10: vec_data_125 = data_d1[79:72];
        7'd11: vec_data_125 = data_d1[87:80];
        7'd12: vec_data_125 = data_d1[95:88];
        7'd13: vec_data_125 = data_d1[103:96];
        7'd14: vec_data_125 = data_d1[111:104];
        7'd15: vec_data_125 = data_d1[119:112];
        7'd16: vec_data_125 = data_d1[127:120];
        7'd17: vec_data_125 = data_d1[135:128];
        7'd18: vec_data_125 = data_d1[143:136];
        7'd19: vec_data_125 = data_d1[151:144];
        7'd20: vec_data_125 = data_d1[159:152];
        7'd21: vec_data_125 = data_d1[167:160];
        7'd22: vec_data_125 = data_d1[175:168];
        7'd23: vec_data_125 = data_d1[183:176];
        7'd24: vec_data_125 = data_d1[191:184];
        7'd25: vec_data_125 = data_d1[199:192];
        7'd26: vec_data_125 = data_d1[207:200];
        7'd27: vec_data_125 = data_d1[215:208];
        7'd28: vec_data_125 = data_d1[223:216];
        7'd29: vec_data_125 = data_d1[231:224];
        7'd30: vec_data_125 = data_d1[239:232];
        7'd31: vec_data_125 = data_d1[247:240];
        7'd32: vec_data_125 = data_d1[255:248];
        7'd33: vec_data_125 = data_d1[263:256];
        7'd34: vec_data_125 = data_d1[271:264];
        7'd35: vec_data_125 = data_d1[279:272];
        7'd36: vec_data_125 = data_d1[287:280];
        7'd37: vec_data_125 = data_d1[295:288];
        7'd38: vec_data_125 = data_d1[303:296];
        7'd39: vec_data_125 = data_d1[311:304];
        7'd40: vec_data_125 = data_d1[319:312];
        7'd41: vec_data_125 = data_d1[327:320];
        7'd42: vec_data_125 = data_d1[335:328];
        7'd43: vec_data_125 = data_d1[343:336];
        7'd44: vec_data_125 = data_d1[351:344];
        7'd45: vec_data_125 = data_d1[359:352];
        7'd46: vec_data_125 = data_d1[367:360];
        7'd47: vec_data_125 = data_d1[375:368];
        7'd48: vec_data_125 = data_d1[383:376];
        7'd49: vec_data_125 = data_d1[391:384];
        7'd50: vec_data_125 = data_d1[399:392];
        7'd51: vec_data_125 = data_d1[407:400];
        7'd52: vec_data_125 = data_d1[415:408];
        7'd53: vec_data_125 = data_d1[423:416];
        7'd54: vec_data_125 = data_d1[431:424];
        7'd55: vec_data_125 = data_d1[439:432];
        7'd56: vec_data_125 = data_d1[447:440];
        7'd57: vec_data_125 = data_d1[455:448];
        7'd58: vec_data_125 = data_d1[463:456];
        7'd59: vec_data_125 = data_d1[471:464];
        7'd60: vec_data_125 = data_d1[479:472];
        7'd61: vec_data_125 = data_d1[487:480];
        7'd62: vec_data_125 = data_d1[495:488];
        7'd63: vec_data_125 = data_d1[503:496];
        7'd64: vec_data_125 = data_d1[511:504];
        7'd65: vec_data_125 = data_d1[519:512];
        7'd66: vec_data_125 = data_d1[527:520];
        7'd67: vec_data_125 = data_d1[535:528];
        7'd68: vec_data_125 = data_d1[543:536];
        7'd69: vec_data_125 = data_d1[551:544];
        7'd70: vec_data_125 = data_d1[559:552];
        7'd71: vec_data_125 = data_d1[567:560];
        7'd72: vec_data_125 = data_d1[575:568];
        7'd73: vec_data_125 = data_d1[583:576];
        7'd74: vec_data_125 = data_d1[591:584];
        7'd75: vec_data_125 = data_d1[599:592];
        7'd76: vec_data_125 = data_d1[607:600];
        7'd77: vec_data_125 = data_d1[615:608];
        7'd78: vec_data_125 = data_d1[623:616];
        7'd79: vec_data_125 = data_d1[631:624];
        7'd80: vec_data_125 = data_d1[639:632];
        7'd81: vec_data_125 = data_d1[647:640];
        7'd82: vec_data_125 = data_d1[655:648];
        7'd83: vec_data_125 = data_d1[663:656];
        7'd84: vec_data_125 = data_d1[671:664];
        7'd85: vec_data_125 = data_d1[679:672];
        7'd86: vec_data_125 = data_d1[687:680];
        7'd87: vec_data_125 = data_d1[695:688];
        7'd88: vec_data_125 = data_d1[703:696];
        7'd89: vec_data_125 = data_d1[711:704];
        7'd90: vec_data_125 = data_d1[719:712];
        7'd91: vec_data_125 = data_d1[727:720];
        7'd92: vec_data_125 = data_d1[735:728];
        7'd93: vec_data_125 = data_d1[743:736];
        7'd94: vec_data_125 = data_d1[751:744];
        7'd95: vec_data_125 = data_d1[759:752];
        7'd96: vec_data_125 = data_d1[767:760];
        7'd97: vec_data_125 = data_d1[775:768];
        7'd98: vec_data_125 = data_d1[783:776];
        7'd99: vec_data_125 = data_d1[791:784];
        7'd100: vec_data_125 = data_d1[799:792];
        7'd101: vec_data_125 = data_d1[807:800];
        7'd102: vec_data_125 = data_d1[815:808];
        7'd103: vec_data_125 = data_d1[823:816];
        7'd104: vec_data_125 = data_d1[831:824];
        7'd105: vec_data_125 = data_d1[839:832];
        7'd106: vec_data_125 = data_d1[847:840];
        7'd107: vec_data_125 = data_d1[855:848];
        7'd108: vec_data_125 = data_d1[863:856];
        7'd109: vec_data_125 = data_d1[871:864];
        7'd110: vec_data_125 = data_d1[879:872];
        7'd111: vec_data_125 = data_d1[887:880];
        7'd112: vec_data_125 = data_d1[895:888];
        7'd113: vec_data_125 = data_d1[903:896];
        7'd114: vec_data_125 = data_d1[911:904];
        7'd115: vec_data_125 = data_d1[919:912];
        7'd116: vec_data_125 = data_d1[927:920];
        7'd117: vec_data_125 = data_d1[935:928];
        7'd118: vec_data_125 = data_d1[943:936];
        7'd119: vec_data_125 = data_d1[951:944];
        7'd120: vec_data_125 = data_d1[959:952];
        7'd121: vec_data_125 = data_d1[967:960];
        7'd122: vec_data_125 = data_d1[975:968];
        7'd123: vec_data_125 = data_d1[983:976];
        7'd124: vec_data_125 = data_d1[991:984];
        7'd125: vec_data_125 = data_d1[999:992];
        7'd126: vec_data_125 = data_d1[1007:1000];
    endcase
end

always @(
  vec_sum_126_d1
  or data_d1
  ) begin
    vec_data_126 = 8'b0;
    case(vec_sum_126_d1)
        7'd1: vec_data_126 = data_d1[7:0];
        7'd2: vec_data_126 = data_d1[15:8];
        7'd3: vec_data_126 = data_d1[23:16];
        7'd4: vec_data_126 = data_d1[31:24];
        7'd5: vec_data_126 = data_d1[39:32];
        7'd6: vec_data_126 = data_d1[47:40];
        7'd7: vec_data_126 = data_d1[55:48];
        7'd8: vec_data_126 = data_d1[63:56];
        7'd9: vec_data_126 = data_d1[71:64];
        7'd10: vec_data_126 = data_d1[79:72];
        7'd11: vec_data_126 = data_d1[87:80];
        7'd12: vec_data_126 = data_d1[95:88];
        7'd13: vec_data_126 = data_d1[103:96];
        7'd14: vec_data_126 = data_d1[111:104];
        7'd15: vec_data_126 = data_d1[119:112];
        7'd16: vec_data_126 = data_d1[127:120];
        7'd17: vec_data_126 = data_d1[135:128];
        7'd18: vec_data_126 = data_d1[143:136];
        7'd19: vec_data_126 = data_d1[151:144];
        7'd20: vec_data_126 = data_d1[159:152];
        7'd21: vec_data_126 = data_d1[167:160];
        7'd22: vec_data_126 = data_d1[175:168];
        7'd23: vec_data_126 = data_d1[183:176];
        7'd24: vec_data_126 = data_d1[191:184];
        7'd25: vec_data_126 = data_d1[199:192];
        7'd26: vec_data_126 = data_d1[207:200];
        7'd27: vec_data_126 = data_d1[215:208];
        7'd28: vec_data_126 = data_d1[223:216];
        7'd29: vec_data_126 = data_d1[231:224];
        7'd30: vec_data_126 = data_d1[239:232];
        7'd31: vec_data_126 = data_d1[247:240];
        7'd32: vec_data_126 = data_d1[255:248];
        7'd33: vec_data_126 = data_d1[263:256];
        7'd34: vec_data_126 = data_d1[271:264];
        7'd35: vec_data_126 = data_d1[279:272];
        7'd36: vec_data_126 = data_d1[287:280];
        7'd37: vec_data_126 = data_d1[295:288];
        7'd38: vec_data_126 = data_d1[303:296];
        7'd39: vec_data_126 = data_d1[311:304];
        7'd40: vec_data_126 = data_d1[319:312];
        7'd41: vec_data_126 = data_d1[327:320];
        7'd42: vec_data_126 = data_d1[335:328];
        7'd43: vec_data_126 = data_d1[343:336];
        7'd44: vec_data_126 = data_d1[351:344];
        7'd45: vec_data_126 = data_d1[359:352];
        7'd46: vec_data_126 = data_d1[367:360];
        7'd47: vec_data_126 = data_d1[375:368];
        7'd48: vec_data_126 = data_d1[383:376];
        7'd49: vec_data_126 = data_d1[391:384];
        7'd50: vec_data_126 = data_d1[399:392];
        7'd51: vec_data_126 = data_d1[407:400];
        7'd52: vec_data_126 = data_d1[415:408];
        7'd53: vec_data_126 = data_d1[423:416];
        7'd54: vec_data_126 = data_d1[431:424];
        7'd55: vec_data_126 = data_d1[439:432];
        7'd56: vec_data_126 = data_d1[447:440];
        7'd57: vec_data_126 = data_d1[455:448];
        7'd58: vec_data_126 = data_d1[463:456];
        7'd59: vec_data_126 = data_d1[471:464];
        7'd60: vec_data_126 = data_d1[479:472];
        7'd61: vec_data_126 = data_d1[487:480];
        7'd62: vec_data_126 = data_d1[495:488];
        7'd63: vec_data_126 = data_d1[503:496];
        7'd64: vec_data_126 = data_d1[511:504];
        7'd65: vec_data_126 = data_d1[519:512];
        7'd66: vec_data_126 = data_d1[527:520];
        7'd67: vec_data_126 = data_d1[535:528];
        7'd68: vec_data_126 = data_d1[543:536];
        7'd69: vec_data_126 = data_d1[551:544];
        7'd70: vec_data_126 = data_d1[559:552];
        7'd71: vec_data_126 = data_d1[567:560];
        7'd72: vec_data_126 = data_d1[575:568];
        7'd73: vec_data_126 = data_d1[583:576];
        7'd74: vec_data_126 = data_d1[591:584];
        7'd75: vec_data_126 = data_d1[599:592];
        7'd76: vec_data_126 = data_d1[607:600];
        7'd77: vec_data_126 = data_d1[615:608];
        7'd78: vec_data_126 = data_d1[623:616];
        7'd79: vec_data_126 = data_d1[631:624];
        7'd80: vec_data_126 = data_d1[639:632];
        7'd81: vec_data_126 = data_d1[647:640];
        7'd82: vec_data_126 = data_d1[655:648];
        7'd83: vec_data_126 = data_d1[663:656];
        7'd84: vec_data_126 = data_d1[671:664];
        7'd85: vec_data_126 = data_d1[679:672];
        7'd86: vec_data_126 = data_d1[687:680];
        7'd87: vec_data_126 = data_d1[695:688];
        7'd88: vec_data_126 = data_d1[703:696];
        7'd89: vec_data_126 = data_d1[711:704];
        7'd90: vec_data_126 = data_d1[719:712];
        7'd91: vec_data_126 = data_d1[727:720];
        7'd92: vec_data_126 = data_d1[735:728];
        7'd93: vec_data_126 = data_d1[743:736];
        7'd94: vec_data_126 = data_d1[751:744];
        7'd95: vec_data_126 = data_d1[759:752];
        7'd96: vec_data_126 = data_d1[767:760];
        7'd97: vec_data_126 = data_d1[775:768];
        7'd98: vec_data_126 = data_d1[783:776];
        7'd99: vec_data_126 = data_d1[791:784];
        7'd100: vec_data_126 = data_d1[799:792];
        7'd101: vec_data_126 = data_d1[807:800];
        7'd102: vec_data_126 = data_d1[815:808];
        7'd103: vec_data_126 = data_d1[823:816];
        7'd104: vec_data_126 = data_d1[831:824];
        7'd105: vec_data_126 = data_d1[839:832];
        7'd106: vec_data_126 = data_d1[847:840];
        7'd107: vec_data_126 = data_d1[855:848];
        7'd108: vec_data_126 = data_d1[863:856];
        7'd109: vec_data_126 = data_d1[871:864];
        7'd110: vec_data_126 = data_d1[879:872];
        7'd111: vec_data_126 = data_d1[887:880];
        7'd112: vec_data_126 = data_d1[895:888];
        7'd113: vec_data_126 = data_d1[903:896];
        7'd114: vec_data_126 = data_d1[911:904];
        7'd115: vec_data_126 = data_d1[919:912];
        7'd116: vec_data_126 = data_d1[927:920];
        7'd117: vec_data_126 = data_d1[935:928];
        7'd118: vec_data_126 = data_d1[943:936];
        7'd119: vec_data_126 = data_d1[951:944];
        7'd120: vec_data_126 = data_d1[959:952];
        7'd121: vec_data_126 = data_d1[967:960];
        7'd122: vec_data_126 = data_d1[975:968];
        7'd123: vec_data_126 = data_d1[983:976];
        7'd124: vec_data_126 = data_d1[991:984];
        7'd125: vec_data_126 = data_d1[999:992];
        7'd126: vec_data_126 = data_d1[1007:1000];
        7'd127: vec_data_126 = data_d1[1015:1008];
    endcase
end

always @(
  vec_sum_127_d1
  or data_d1
  ) begin
    vec_data_127 = 8'b0;
    case(vec_sum_127_d1)
        8'd1: vec_data_127 = data_d1[7:0];
        8'd2: vec_data_127 = data_d1[15:8];
        8'd3: vec_data_127 = data_d1[23:16];
        8'd4: vec_data_127 = data_d1[31:24];
        8'd5: vec_data_127 = data_d1[39:32];
        8'd6: vec_data_127 = data_d1[47:40];
        8'd7: vec_data_127 = data_d1[55:48];
        8'd8: vec_data_127 = data_d1[63:56];
        8'd9: vec_data_127 = data_d1[71:64];
        8'd10: vec_data_127 = data_d1[79:72];
        8'd11: vec_data_127 = data_d1[87:80];
        8'd12: vec_data_127 = data_d1[95:88];
        8'd13: vec_data_127 = data_d1[103:96];
        8'd14: vec_data_127 = data_d1[111:104];
        8'd15: vec_data_127 = data_d1[119:112];
        8'd16: vec_data_127 = data_d1[127:120];
        8'd17: vec_data_127 = data_d1[135:128];
        8'd18: vec_data_127 = data_d1[143:136];
        8'd19: vec_data_127 = data_d1[151:144];
        8'd20: vec_data_127 = data_d1[159:152];
        8'd21: vec_data_127 = data_d1[167:160];
        8'd22: vec_data_127 = data_d1[175:168];
        8'd23: vec_data_127 = data_d1[183:176];
        8'd24: vec_data_127 = data_d1[191:184];
        8'd25: vec_data_127 = data_d1[199:192];
        8'd26: vec_data_127 = data_d1[207:200];
        8'd27: vec_data_127 = data_d1[215:208];
        8'd28: vec_data_127 = data_d1[223:216];
        8'd29: vec_data_127 = data_d1[231:224];
        8'd30: vec_data_127 = data_d1[239:232];
        8'd31: vec_data_127 = data_d1[247:240];
        8'd32: vec_data_127 = data_d1[255:248];
        8'd33: vec_data_127 = data_d1[263:256];
        8'd34: vec_data_127 = data_d1[271:264];
        8'd35: vec_data_127 = data_d1[279:272];
        8'd36: vec_data_127 = data_d1[287:280];
        8'd37: vec_data_127 = data_d1[295:288];
        8'd38: vec_data_127 = data_d1[303:296];
        8'd39: vec_data_127 = data_d1[311:304];
        8'd40: vec_data_127 = data_d1[319:312];
        8'd41: vec_data_127 = data_d1[327:320];
        8'd42: vec_data_127 = data_d1[335:328];
        8'd43: vec_data_127 = data_d1[343:336];
        8'd44: vec_data_127 = data_d1[351:344];
        8'd45: vec_data_127 = data_d1[359:352];
        8'd46: vec_data_127 = data_d1[367:360];
        8'd47: vec_data_127 = data_d1[375:368];
        8'd48: vec_data_127 = data_d1[383:376];
        8'd49: vec_data_127 = data_d1[391:384];
        8'd50: vec_data_127 = data_d1[399:392];
        8'd51: vec_data_127 = data_d1[407:400];
        8'd52: vec_data_127 = data_d1[415:408];
        8'd53: vec_data_127 = data_d1[423:416];
        8'd54: vec_data_127 = data_d1[431:424];
        8'd55: vec_data_127 = data_d1[439:432];
        8'd56: vec_data_127 = data_d1[447:440];
        8'd57: vec_data_127 = data_d1[455:448];
        8'd58: vec_data_127 = data_d1[463:456];
        8'd59: vec_data_127 = data_d1[471:464];
        8'd60: vec_data_127 = data_d1[479:472];
        8'd61: vec_data_127 = data_d1[487:480];
        8'd62: vec_data_127 = data_d1[495:488];
        8'd63: vec_data_127 = data_d1[503:496];
        8'd64: vec_data_127 = data_d1[511:504];
        8'd65: vec_data_127 = data_d1[519:512];
        8'd66: vec_data_127 = data_d1[527:520];
        8'd67: vec_data_127 = data_d1[535:528];
        8'd68: vec_data_127 = data_d1[543:536];
        8'd69: vec_data_127 = data_d1[551:544];
        8'd70: vec_data_127 = data_d1[559:552];
        8'd71: vec_data_127 = data_d1[567:560];
        8'd72: vec_data_127 = data_d1[575:568];
        8'd73: vec_data_127 = data_d1[583:576];
        8'd74: vec_data_127 = data_d1[591:584];
        8'd75: vec_data_127 = data_d1[599:592];
        8'd76: vec_data_127 = data_d1[607:600];
        8'd77: vec_data_127 = data_d1[615:608];
        8'd78: vec_data_127 = data_d1[623:616];
        8'd79: vec_data_127 = data_d1[631:624];
        8'd80: vec_data_127 = data_d1[639:632];
        8'd81: vec_data_127 = data_d1[647:640];
        8'd82: vec_data_127 = data_d1[655:648];
        8'd83: vec_data_127 = data_d1[663:656];
        8'd84: vec_data_127 = data_d1[671:664];
        8'd85: vec_data_127 = data_d1[679:672];
        8'd86: vec_data_127 = data_d1[687:680];
        8'd87: vec_data_127 = data_d1[695:688];
        8'd88: vec_data_127 = data_d1[703:696];
        8'd89: vec_data_127 = data_d1[711:704];
        8'd90: vec_data_127 = data_d1[719:712];
        8'd91: vec_data_127 = data_d1[727:720];
        8'd92: vec_data_127 = data_d1[735:728];
        8'd93: vec_data_127 = data_d1[743:736];
        8'd94: vec_data_127 = data_d1[751:744];
        8'd95: vec_data_127 = data_d1[759:752];
        8'd96: vec_data_127 = data_d1[767:760];
        8'd97: vec_data_127 = data_d1[775:768];
        8'd98: vec_data_127 = data_d1[783:776];
        8'd99: vec_data_127 = data_d1[791:784];
        8'd100: vec_data_127 = data_d1[799:792];
        8'd101: vec_data_127 = data_d1[807:800];
        8'd102: vec_data_127 = data_d1[815:808];
        8'd103: vec_data_127 = data_d1[823:816];
        8'd104: vec_data_127 = data_d1[831:824];
        8'd105: vec_data_127 = data_d1[839:832];
        8'd106: vec_data_127 = data_d1[847:840];
        8'd107: vec_data_127 = data_d1[855:848];
        8'd108: vec_data_127 = data_d1[863:856];
        8'd109: vec_data_127 = data_d1[871:864];
        8'd110: vec_data_127 = data_d1[879:872];
        8'd111: vec_data_127 = data_d1[887:880];
        8'd112: vec_data_127 = data_d1[895:888];
        8'd113: vec_data_127 = data_d1[903:896];
        8'd114: vec_data_127 = data_d1[911:904];
        8'd115: vec_data_127 = data_d1[919:912];
        8'd116: vec_data_127 = data_d1[927:920];
        8'd117: vec_data_127 = data_d1[935:928];
        8'd118: vec_data_127 = data_d1[943:936];
        8'd119: vec_data_127 = data_d1[951:944];
        8'd120: vec_data_127 = data_d1[959:952];
        8'd121: vec_data_127 = data_d1[967:960];
        8'd122: vec_data_127 = data_d1[975:968];
        8'd123: vec_data_127 = data_d1[983:976];
        8'd124: vec_data_127 = data_d1[991:984];
        8'd125: vec_data_127 = data_d1[999:992];
        8'd126: vec_data_127 = data_d1[1007:1000];
        8'd127: vec_data_127 = data_d1[1015:1008];
        8'd128: vec_data_127 = data_d1[1023:1016];
    endcase
end



////////////////////////////////// phase II: registers and assertion //////////////////////////////////
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    valid_d2 <= 1'b0;
  end else begin
  valid_d2 <= valid_d1;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    sel_d2 <= sel_d1;
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    sel_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_000_d2 <= (vec_data_000 & {8{mask_d1[0]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_000_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_001_d2 <= (vec_data_001 & {8{mask_d1[1]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_001_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_002_d2 <= (vec_data_002 & {8{mask_d1[2]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_002_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_003_d2 <= (vec_data_003 & {8{mask_d1[3]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_003_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_004_d2 <= (vec_data_004 & {8{mask_d1[4]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_004_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_005_d2 <= (vec_data_005 & {8{mask_d1[5]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_005_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_006_d2 <= (vec_data_006 & {8{mask_d1[6]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_006_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_007_d2 <= (vec_data_007 & {8{mask_d1[7]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_007_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_008_d2 <= (vec_data_008 & {8{mask_d1[8]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_008_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_009_d2 <= (vec_data_009 & {8{mask_d1[9]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_009_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_010_d2 <= (vec_data_010 & {8{mask_d1[10]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_010_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_011_d2 <= (vec_data_011 & {8{mask_d1[11]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_011_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_012_d2 <= (vec_data_012 & {8{mask_d1[12]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_012_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_013_d2 <= (vec_data_013 & {8{mask_d1[13]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_013_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_014_d2 <= (vec_data_014 & {8{mask_d1[14]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_014_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_015_d2 <= (vec_data_015 & {8{mask_d1[15]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_015_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_016_d2 <= (vec_data_016 & {8{mask_d1[16]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_016_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_017_d2 <= (vec_data_017 & {8{mask_d1[17]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_017_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_018_d2 <= (vec_data_018 & {8{mask_d1[18]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_018_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_019_d2 <= (vec_data_019 & {8{mask_d1[19]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_019_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_020_d2 <= (vec_data_020 & {8{mask_d1[20]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_020_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_021_d2 <= (vec_data_021 & {8{mask_d1[21]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_021_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_022_d2 <= (vec_data_022 & {8{mask_d1[22]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_022_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_023_d2 <= (vec_data_023 & {8{mask_d1[23]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_023_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_024_d2 <= (vec_data_024 & {8{mask_d1[24]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_024_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_025_d2 <= (vec_data_025 & {8{mask_d1[25]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_025_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_026_d2 <= (vec_data_026 & {8{mask_d1[26]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_026_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_027_d2 <= (vec_data_027 & {8{mask_d1[27]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_027_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_028_d2 <= (vec_data_028 & {8{mask_d1[28]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_028_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_029_d2 <= (vec_data_029 & {8{mask_d1[29]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_029_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_030_d2 <= (vec_data_030 & {8{mask_d1[30]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_030_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_031_d2 <= (vec_data_031 & {8{mask_d1[31]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_031_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_032_d2 <= (vec_data_032 & {8{mask_d1[32]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_032_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_033_d2 <= (vec_data_033 & {8{mask_d1[33]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_033_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_034_d2 <= (vec_data_034 & {8{mask_d1[34]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_034_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_035_d2 <= (vec_data_035 & {8{mask_d1[35]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_035_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_036_d2 <= (vec_data_036 & {8{mask_d1[36]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_036_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_037_d2 <= (vec_data_037 & {8{mask_d1[37]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_037_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_038_d2 <= (vec_data_038 & {8{mask_d1[38]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_038_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_039_d2 <= (vec_data_039 & {8{mask_d1[39]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_039_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_040_d2 <= (vec_data_040 & {8{mask_d1[40]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_040_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_041_d2 <= (vec_data_041 & {8{mask_d1[41]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_041_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_042_d2 <= (vec_data_042 & {8{mask_d1[42]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_042_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_043_d2 <= (vec_data_043 & {8{mask_d1[43]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_043_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_044_d2 <= (vec_data_044 & {8{mask_d1[44]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_044_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_045_d2 <= (vec_data_045 & {8{mask_d1[45]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_045_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_046_d2 <= (vec_data_046 & {8{mask_d1[46]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_046_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_047_d2 <= (vec_data_047 & {8{mask_d1[47]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_047_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_048_d2 <= (vec_data_048 & {8{mask_d1[48]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_048_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_049_d2 <= (vec_data_049 & {8{mask_d1[49]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_049_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_050_d2 <= (vec_data_050 & {8{mask_d1[50]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_050_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_051_d2 <= (vec_data_051 & {8{mask_d1[51]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_051_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_052_d2 <= (vec_data_052 & {8{mask_d1[52]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_052_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_053_d2 <= (vec_data_053 & {8{mask_d1[53]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_053_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_054_d2 <= (vec_data_054 & {8{mask_d1[54]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_054_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_055_d2 <= (vec_data_055 & {8{mask_d1[55]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_055_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_056_d2 <= (vec_data_056 & {8{mask_d1[56]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_056_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_057_d2 <= (vec_data_057 & {8{mask_d1[57]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_057_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_058_d2 <= (vec_data_058 & {8{mask_d1[58]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_058_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_059_d2 <= (vec_data_059 & {8{mask_d1[59]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_059_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_060_d2 <= (vec_data_060 & {8{mask_d1[60]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_060_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_061_d2 <= (vec_data_061 & {8{mask_d1[61]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_061_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_062_d2 <= (vec_data_062 & {8{mask_d1[62]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_062_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_063_d2 <= (vec_data_063 & {8{mask_d1[63]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_063_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_064_d2 <= (vec_data_064 & {8{mask_d1[64]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_064_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_065_d2 <= (vec_data_065 & {8{mask_d1[65]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_065_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_066_d2 <= (vec_data_066 & {8{mask_d1[66]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_066_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_067_d2 <= (vec_data_067 & {8{mask_d1[67]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_067_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_068_d2 <= (vec_data_068 & {8{mask_d1[68]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_068_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_069_d2 <= (vec_data_069 & {8{mask_d1[69]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_069_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_070_d2 <= (vec_data_070 & {8{mask_d1[70]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_070_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_071_d2 <= (vec_data_071 & {8{mask_d1[71]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_071_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_072_d2 <= (vec_data_072 & {8{mask_d1[72]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_072_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_073_d2 <= (vec_data_073 & {8{mask_d1[73]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_073_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_074_d2 <= (vec_data_074 & {8{mask_d1[74]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_074_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_075_d2 <= (vec_data_075 & {8{mask_d1[75]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_075_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_076_d2 <= (vec_data_076 & {8{mask_d1[76]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_076_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_077_d2 <= (vec_data_077 & {8{mask_d1[77]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_077_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_078_d2 <= (vec_data_078 & {8{mask_d1[78]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_078_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_079_d2 <= (vec_data_079 & {8{mask_d1[79]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_079_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_080_d2 <= (vec_data_080 & {8{mask_d1[80]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_080_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_081_d2 <= (vec_data_081 & {8{mask_d1[81]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_081_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_082_d2 <= (vec_data_082 & {8{mask_d1[82]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_082_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_083_d2 <= (vec_data_083 & {8{mask_d1[83]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_083_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_084_d2 <= (vec_data_084 & {8{mask_d1[84]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_084_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_085_d2 <= (vec_data_085 & {8{mask_d1[85]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_085_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_086_d2 <= (vec_data_086 & {8{mask_d1[86]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_086_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_087_d2 <= (vec_data_087 & {8{mask_d1[87]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_087_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_088_d2 <= (vec_data_088 & {8{mask_d1[88]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_088_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_089_d2 <= (vec_data_089 & {8{mask_d1[89]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_089_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_090_d2 <= (vec_data_090 & {8{mask_d1[90]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_090_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_091_d2 <= (vec_data_091 & {8{mask_d1[91]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_091_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_092_d2 <= (vec_data_092 & {8{mask_d1[92]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_092_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_093_d2 <= (vec_data_093 & {8{mask_d1[93]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_093_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_094_d2 <= (vec_data_094 & {8{mask_d1[94]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_094_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_095_d2 <= (vec_data_095 & {8{mask_d1[95]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_095_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_096_d2 <= (vec_data_096 & {8{mask_d1[96]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_096_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_097_d2 <= (vec_data_097 & {8{mask_d1[97]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_097_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_098_d2 <= (vec_data_098 & {8{mask_d1[98]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_098_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_099_d2 <= (vec_data_099 & {8{mask_d1[99]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_099_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_100_d2 <= (vec_data_100 & {8{mask_d1[100]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_100_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_101_d2 <= (vec_data_101 & {8{mask_d1[101]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_101_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_102_d2 <= (vec_data_102 & {8{mask_d1[102]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_102_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_103_d2 <= (vec_data_103 & {8{mask_d1[103]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_103_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_104_d2 <= (vec_data_104 & {8{mask_d1[104]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_104_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_105_d2 <= (vec_data_105 & {8{mask_d1[105]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_105_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_106_d2 <= (vec_data_106 & {8{mask_d1[106]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_106_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_107_d2 <= (vec_data_107 & {8{mask_d1[107]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_107_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_108_d2 <= (vec_data_108 & {8{mask_d1[108]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_108_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_109_d2 <= (vec_data_109 & {8{mask_d1[109]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_109_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_110_d2 <= (vec_data_110 & {8{mask_d1[110]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_110_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_111_d2 <= (vec_data_111 & {8{mask_d1[111]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_111_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_112_d2 <= (vec_data_112 & {8{mask_d1[112]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_112_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_113_d2 <= (vec_data_113 & {8{mask_d1[113]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_113_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_114_d2 <= (vec_data_114 & {8{mask_d1[114]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_114_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_115_d2 <= (vec_data_115 & {8{mask_d1[115]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_115_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_116_d2 <= (vec_data_116 & {8{mask_d1[116]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_116_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_117_d2 <= (vec_data_117 & {8{mask_d1[117]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_117_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_118_d2 <= (vec_data_118 & {8{mask_d1[118]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_118_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_119_d2 <= (vec_data_119 & {8{mask_d1[119]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_119_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_120_d2 <= (vec_data_120 & {8{mask_d1[120]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_120_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_121_d2 <= (vec_data_121 & {8{mask_d1[121]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_121_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_122_d2 <= (vec_data_122 & {8{mask_d1[122]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_122_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_123_d2 <= (vec_data_123 & {8{mask_d1[123]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_123_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_124_d2 <= (vec_data_124 & {8{mask_d1[124]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_124_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_125_d2 <= (vec_data_125 & {8{mask_d1[125]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_125_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_126_d2 <= (vec_data_126 & {8{mask_d1[126]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_126_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d1) == 1'b1) begin
    vec_data_127_d2 <= (vec_data_127 & {8{mask_d1[127]}});
  // VCS coverage off
  end else if ((valid_d1) == 1'b0) begin
  end else begin
    vec_data_127_d2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_000_d1 is out of range! ")      zzz_assert_never_1x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_000_d1 > 1'd1))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_001_d1 is out of range! ")      zzz_assert_never_2x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_001_d1 > 2'd2))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_002_d1 is out of range! ")      zzz_assert_never_3x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_002_d1 > 2'd3))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_003_d1 is out of range! ")      zzz_assert_never_4x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_003_d1 > 3'd4))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_004_d1 is out of range! ")      zzz_assert_never_5x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_004_d1 > 3'd5))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_005_d1 is out of range! ")      zzz_assert_never_6x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_005_d1 > 3'd6))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_006_d1 is out of range! ")      zzz_assert_never_7x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_006_d1 > 3'd7))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_007_d1 is out of range! ")      zzz_assert_never_8x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_007_d1 > 4'd8))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_008_d1 is out of range! ")      zzz_assert_never_9x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_008_d1 > 4'd9))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_009_d1 is out of range! ")      zzz_assert_never_10x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_009_d1 > 4'd10))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_010_d1 is out of range! ")      zzz_assert_never_11x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_010_d1 > 4'd11))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_011_d1 is out of range! ")      zzz_assert_never_12x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_011_d1 > 4'd12))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_012_d1 is out of range! ")      zzz_assert_never_13x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_012_d1 > 4'd13))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_013_d1 is out of range! ")      zzz_assert_never_14x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_013_d1 > 4'd14))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_014_d1 is out of range! ")      zzz_assert_never_15x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_014_d1 > 4'd15))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_015_d1 is out of range! ")      zzz_assert_never_16x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_015_d1 > 5'd16))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_016_d1 is out of range! ")      zzz_assert_never_17x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_016_d1 > 5'd17))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_017_d1 is out of range! ")      zzz_assert_never_18x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_017_d1 > 5'd18))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_018_d1 is out of range! ")      zzz_assert_never_19x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_018_d1 > 5'd19))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_019_d1 is out of range! ")      zzz_assert_never_20x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_019_d1 > 5'd20))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_020_d1 is out of range! ")      zzz_assert_never_21x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_020_d1 > 5'd21))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_021_d1 is out of range! ")      zzz_assert_never_22x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_021_d1 > 5'd22))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_022_d1 is out of range! ")      zzz_assert_never_23x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_022_d1 > 5'd23))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_023_d1 is out of range! ")      zzz_assert_never_24x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_023_d1 > 5'd24))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_024_d1 is out of range! ")      zzz_assert_never_25x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_024_d1 > 5'd25))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_025_d1 is out of range! ")      zzz_assert_never_26x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_025_d1 > 5'd26))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_026_d1 is out of range! ")      zzz_assert_never_27x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_026_d1 > 5'd27))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_027_d1 is out of range! ")      zzz_assert_never_28x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_027_d1 > 5'd28))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_028_d1 is out of range! ")      zzz_assert_never_29x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_028_d1 > 5'd29))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_029_d1 is out of range! ")      zzz_assert_never_30x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_029_d1 > 5'd30))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_030_d1 is out of range! ")      zzz_assert_never_31x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_030_d1 > 5'd31))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_031_d1 is out of range! ")      zzz_assert_never_32x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_031_d1 > 6'd32))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_032_d1 is out of range! ")      zzz_assert_never_33x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_032_d1 > 6'd33))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_033_d1 is out of range! ")      zzz_assert_never_34x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_033_d1 > 6'd34))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_034_d1 is out of range! ")      zzz_assert_never_35x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_034_d1 > 6'd35))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_035_d1 is out of range! ")      zzz_assert_never_36x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_035_d1 > 6'd36))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_036_d1 is out of range! ")      zzz_assert_never_37x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_036_d1 > 6'd37))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_037_d1 is out of range! ")      zzz_assert_never_38x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_037_d1 > 6'd38))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_038_d1 is out of range! ")      zzz_assert_never_39x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_038_d1 > 6'd39))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_039_d1 is out of range! ")      zzz_assert_never_40x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_039_d1 > 6'd40))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_040_d1 is out of range! ")      zzz_assert_never_41x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_040_d1 > 6'd41))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_041_d1 is out of range! ")      zzz_assert_never_42x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_041_d1 > 6'd42))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_042_d1 is out of range! ")      zzz_assert_never_43x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_042_d1 > 6'd43))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_043_d1 is out of range! ")      zzz_assert_never_44x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_043_d1 > 6'd44))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_044_d1 is out of range! ")      zzz_assert_never_45x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_044_d1 > 6'd45))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_045_d1 is out of range! ")      zzz_assert_never_46x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_045_d1 > 6'd46))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_046_d1 is out of range! ")      zzz_assert_never_47x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_046_d1 > 6'd47))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_047_d1 is out of range! ")      zzz_assert_never_48x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_047_d1 > 6'd48))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_048_d1 is out of range! ")      zzz_assert_never_49x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_048_d1 > 6'd49))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_049_d1 is out of range! ")      zzz_assert_never_50x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_049_d1 > 6'd50))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_050_d1 is out of range! ")      zzz_assert_never_51x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_050_d1 > 6'd51))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_051_d1 is out of range! ")      zzz_assert_never_52x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_051_d1 > 6'd52))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_052_d1 is out of range! ")      zzz_assert_never_53x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_052_d1 > 6'd53))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_053_d1 is out of range! ")      zzz_assert_never_54x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_053_d1 > 6'd54))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_054_d1 is out of range! ")      zzz_assert_never_55x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_054_d1 > 6'd55))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_055_d1 is out of range! ")      zzz_assert_never_56x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_055_d1 > 6'd56))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_056_d1 is out of range! ")      zzz_assert_never_57x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_056_d1 > 6'd57))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_057_d1 is out of range! ")      zzz_assert_never_58x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_057_d1 > 6'd58))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_058_d1 is out of range! ")      zzz_assert_never_59x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_058_d1 > 6'd59))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_059_d1 is out of range! ")      zzz_assert_never_60x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_059_d1 > 6'd60))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_060_d1 is out of range! ")      zzz_assert_never_61x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_060_d1 > 6'd61))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_061_d1 is out of range! ")      zzz_assert_never_62x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_061_d1 > 6'd62))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_062_d1 is out of range! ")      zzz_assert_never_63x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_062_d1 > 6'd63))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_063_d1 is out of range! ")      zzz_assert_never_64x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_063_d1 > 7'd64))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_064_d1 is out of range! ")      zzz_assert_never_65x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_064_d1 > 7'd65))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_065_d1 is out of range! ")      zzz_assert_never_66x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_065_d1 > 7'd66))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_066_d1 is out of range! ")      zzz_assert_never_67x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_066_d1 > 7'd67))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_067_d1 is out of range! ")      zzz_assert_never_68x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_067_d1 > 7'd68))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_068_d1 is out of range! ")      zzz_assert_never_69x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_068_d1 > 7'd69))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_069_d1 is out of range! ")      zzz_assert_never_70x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_069_d1 > 7'd70))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_070_d1 is out of range! ")      zzz_assert_never_71x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_070_d1 > 7'd71))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_071_d1 is out of range! ")      zzz_assert_never_72x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_071_d1 > 7'd72))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_072_d1 is out of range! ")      zzz_assert_never_73x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_072_d1 > 7'd73))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_073_d1 is out of range! ")      zzz_assert_never_74x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_073_d1 > 7'd74))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_074_d1 is out of range! ")      zzz_assert_never_75x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_074_d1 > 7'd75))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_075_d1 is out of range! ")      zzz_assert_never_76x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_075_d1 > 7'd76))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_076_d1 is out of range! ")      zzz_assert_never_77x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_076_d1 > 7'd77))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_077_d1 is out of range! ")      zzz_assert_never_78x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_077_d1 > 7'd78))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_078_d1 is out of range! ")      zzz_assert_never_79x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_078_d1 > 7'd79))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_079_d1 is out of range! ")      zzz_assert_never_80x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_079_d1 > 7'd80))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_080_d1 is out of range! ")      zzz_assert_never_81x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_080_d1 > 7'd81))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_081_d1 is out of range! ")      zzz_assert_never_82x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_081_d1 > 7'd82))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_082_d1 is out of range! ")      zzz_assert_never_83x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_082_d1 > 7'd83))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_083_d1 is out of range! ")      zzz_assert_never_84x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_083_d1 > 7'd84))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_084_d1 is out of range! ")      zzz_assert_never_85x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_084_d1 > 7'd85))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_085_d1 is out of range! ")      zzz_assert_never_86x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_085_d1 > 7'd86))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_086_d1 is out of range! ")      zzz_assert_never_87x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_086_d1 > 7'd87))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_087_d1 is out of range! ")      zzz_assert_never_88x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_087_d1 > 7'd88))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_088_d1 is out of range! ")      zzz_assert_never_89x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_088_d1 > 7'd89))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_089_d1 is out of range! ")      zzz_assert_never_90x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_089_d1 > 7'd90))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_090_d1 is out of range! ")      zzz_assert_never_91x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_090_d1 > 7'd91))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_091_d1 is out of range! ")      zzz_assert_never_92x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_091_d1 > 7'd92))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_092_d1 is out of range! ")      zzz_assert_never_93x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_092_d1 > 7'd93))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_093_d1 is out of range! ")      zzz_assert_never_94x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_093_d1 > 7'd94))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_094_d1 is out of range! ")      zzz_assert_never_95x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_094_d1 > 7'd95))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_095_d1 is out of range! ")      zzz_assert_never_96x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_095_d1 > 7'd96))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_096_d1 is out of range! ")      zzz_assert_never_97x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_096_d1 > 7'd97))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_097_d1 is out of range! ")      zzz_assert_never_98x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_097_d1 > 7'd98))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_098_d1 is out of range! ")      zzz_assert_never_99x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_098_d1 > 7'd99))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_099_d1 is out of range! ")      zzz_assert_never_100x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_099_d1 > 7'd100))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_100_d1 is out of range! ")      zzz_assert_never_101x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_100_d1 > 7'd101))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_101_d1 is out of range! ")      zzz_assert_never_102x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_101_d1 > 7'd102))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_102_d1 is out of range! ")      zzz_assert_never_103x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_102_d1 > 7'd103))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_103_d1 is out of range! ")      zzz_assert_never_104x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_103_d1 > 7'd104))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_104_d1 is out of range! ")      zzz_assert_never_105x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_104_d1 > 7'd105))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_105_d1 is out of range! ")      zzz_assert_never_106x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_105_d1 > 7'd106))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_106_d1 is out of range! ")      zzz_assert_never_107x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_106_d1 > 7'd107))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_107_d1 is out of range! ")      zzz_assert_never_108x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_107_d1 > 7'd108))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_108_d1 is out of range! ")      zzz_assert_never_109x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_108_d1 > 7'd109))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_109_d1 is out of range! ")      zzz_assert_never_110x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_109_d1 > 7'd110))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_110_d1 is out of range! ")      zzz_assert_never_111x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_110_d1 > 7'd111))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_111_d1 is out of range! ")      zzz_assert_never_112x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_111_d1 > 7'd112))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_112_d1 is out of range! ")      zzz_assert_never_113x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_112_d1 > 7'd113))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_113_d1 is out of range! ")      zzz_assert_never_114x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_113_d1 > 7'd114))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_114_d1 is out of range! ")      zzz_assert_never_115x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_114_d1 > 7'd115))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_115_d1 is out of range! ")      zzz_assert_never_116x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_115_d1 > 7'd116))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_116_d1 is out of range! ")      zzz_assert_never_117x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_116_d1 > 7'd117))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_117_d1 is out of range! ")      zzz_assert_never_118x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_117_d1 > 7'd118))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_118_d1 is out of range! ")      zzz_assert_never_119x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_118_d1 > 7'd119))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_119_d1 is out of range! ")      zzz_assert_never_120x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_119_d1 > 7'd120))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_120_d1 is out of range! ")      zzz_assert_never_121x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_120_d1 > 7'd121))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_121_d1 is out of range! ")      zzz_assert_never_122x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_121_d1 > 7'd122))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_122_d1 is out of range! ")      zzz_assert_never_123x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_122_d1 > 7'd123))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_123_d1 is out of range! ")      zzz_assert_never_124x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_123_d1 > 7'd124))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_124_d1 is out of range! ")      zzz_assert_never_125x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_124_d1 > 7'd125))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_125_d1 is out of range! ")      zzz_assert_never_126x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_125_d1 > 7'd126))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_126_d1 is out of range! ")      zzz_assert_never_127x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_126_d1 > 7'd127))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error!  vec_sum_127_d1 is out of range! ")      zzz_assert_never_128x (nvdla_core_clk, `ASSERT_RESET, (valid_d1 && (vec_sum_127_d1 > 8'd128))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
////////////////////////////////// phase III: registers //////////////////////////////////
always @(
  vec_data_000_d2
  or vec_data_001_d2
  or vec_data_002_d2
  or vec_data_003_d2
  or vec_data_004_d2
  or vec_data_005_d2
  or vec_data_006_d2
  or vec_data_007_d2
  or vec_data_008_d2
  or vec_data_009_d2
  or vec_data_010_d2
  or vec_data_011_d2
  or vec_data_012_d2
  or vec_data_013_d2
  or vec_data_014_d2
  or vec_data_015_d2
  or vec_data_016_d2
  or vec_data_017_d2
  or vec_data_018_d2
  or vec_data_019_d2
  or vec_data_020_d2
  or vec_data_021_d2
  or vec_data_022_d2
  or vec_data_023_d2
  or vec_data_024_d2
  or vec_data_025_d2
  or vec_data_026_d2
  or vec_data_027_d2
  or vec_data_028_d2
  or vec_data_029_d2
  or vec_data_030_d2
  or vec_data_031_d2
  or vec_data_032_d2
  or vec_data_033_d2
  or vec_data_034_d2
  or vec_data_035_d2
  or vec_data_036_d2
  or vec_data_037_d2
  or vec_data_038_d2
  or vec_data_039_d2
  or vec_data_040_d2
  or vec_data_041_d2
  or vec_data_042_d2
  or vec_data_043_d2
  or vec_data_044_d2
  or vec_data_045_d2
  or vec_data_046_d2
  or vec_data_047_d2
  or vec_data_048_d2
  or vec_data_049_d2
  or vec_data_050_d2
  or vec_data_051_d2
  or vec_data_052_d2
  or vec_data_053_d2
  or vec_data_054_d2
  or vec_data_055_d2
  or vec_data_056_d2
  or vec_data_057_d2
  or vec_data_058_d2
  or vec_data_059_d2
  or vec_data_060_d2
  or vec_data_061_d2
  or vec_data_062_d2
  or vec_data_063_d2
  or vec_data_064_d2
  or vec_data_065_d2
  or vec_data_066_d2
  or vec_data_067_d2
  or vec_data_068_d2
  or vec_data_069_d2
  or vec_data_070_d2
  or vec_data_071_d2
  or vec_data_072_d2
  or vec_data_073_d2
  or vec_data_074_d2
  or vec_data_075_d2
  or vec_data_076_d2
  or vec_data_077_d2
  or vec_data_078_d2
  or vec_data_079_d2
  or vec_data_080_d2
  or vec_data_081_d2
  or vec_data_082_d2
  or vec_data_083_d2
  or vec_data_084_d2
  or vec_data_085_d2
  or vec_data_086_d2
  or vec_data_087_d2
  or vec_data_088_d2
  or vec_data_089_d2
  or vec_data_090_d2
  or vec_data_091_d2
  or vec_data_092_d2
  or vec_data_093_d2
  or vec_data_094_d2
  or vec_data_095_d2
  or vec_data_096_d2
  or vec_data_097_d2
  or vec_data_098_d2
  or vec_data_099_d2
  or vec_data_100_d2
  or vec_data_101_d2
  or vec_data_102_d2
  or vec_data_103_d2
  or vec_data_104_d2
  or vec_data_105_d2
  or vec_data_106_d2
  or vec_data_107_d2
  or vec_data_108_d2
  or vec_data_109_d2
  or vec_data_110_d2
  or vec_data_111_d2
  or vec_data_112_d2
  or vec_data_113_d2
  or vec_data_114_d2
  or vec_data_115_d2
  or vec_data_116_d2
  or vec_data_117_d2
  or vec_data_118_d2
  or vec_data_119_d2
  or vec_data_120_d2
  or vec_data_121_d2
  or vec_data_122_d2
  or vec_data_123_d2
  or vec_data_124_d2
  or vec_data_125_d2
  or vec_data_126_d2
  or vec_data_127_d2
  ) begin
    mask_d2_int8_w[0] = (|vec_data_000_d2);
    mask_d2_int8_w[1] = (|vec_data_001_d2);
    mask_d2_int8_w[2] = (|vec_data_002_d2);
    mask_d2_int8_w[3] = (|vec_data_003_d2);
    mask_d2_int8_w[4] = (|vec_data_004_d2);
    mask_d2_int8_w[5] = (|vec_data_005_d2);
    mask_d2_int8_w[6] = (|vec_data_006_d2);
    mask_d2_int8_w[7] = (|vec_data_007_d2);
    mask_d2_int8_w[8] = (|vec_data_008_d2);
    mask_d2_int8_w[9] = (|vec_data_009_d2);
    mask_d2_int8_w[10] = (|vec_data_010_d2);
    mask_d2_int8_w[11] = (|vec_data_011_d2);
    mask_d2_int8_w[12] = (|vec_data_012_d2);
    mask_d2_int8_w[13] = (|vec_data_013_d2);
    mask_d2_int8_w[14] = (|vec_data_014_d2);
    mask_d2_int8_w[15] = (|vec_data_015_d2);
    mask_d2_int8_w[16] = (|vec_data_016_d2);
    mask_d2_int8_w[17] = (|vec_data_017_d2);
    mask_d2_int8_w[18] = (|vec_data_018_d2);
    mask_d2_int8_w[19] = (|vec_data_019_d2);
    mask_d2_int8_w[20] = (|vec_data_020_d2);
    mask_d2_int8_w[21] = (|vec_data_021_d2);
    mask_d2_int8_w[22] = (|vec_data_022_d2);
    mask_d2_int8_w[23] = (|vec_data_023_d2);
    mask_d2_int8_w[24] = (|vec_data_024_d2);
    mask_d2_int8_w[25] = (|vec_data_025_d2);
    mask_d2_int8_w[26] = (|vec_data_026_d2);
    mask_d2_int8_w[27] = (|vec_data_027_d2);
    mask_d2_int8_w[28] = (|vec_data_028_d2);
    mask_d2_int8_w[29] = (|vec_data_029_d2);
    mask_d2_int8_w[30] = (|vec_data_030_d2);
    mask_d2_int8_w[31] = (|vec_data_031_d2);
    mask_d2_int8_w[32] = (|vec_data_032_d2);
    mask_d2_int8_w[33] = (|vec_data_033_d2);
    mask_d2_int8_w[34] = (|vec_data_034_d2);
    mask_d2_int8_w[35] = (|vec_data_035_d2);
    mask_d2_int8_w[36] = (|vec_data_036_d2);
    mask_d2_int8_w[37] = (|vec_data_037_d2);
    mask_d2_int8_w[38] = (|vec_data_038_d2);
    mask_d2_int8_w[39] = (|vec_data_039_d2);
    mask_d2_int8_w[40] = (|vec_data_040_d2);
    mask_d2_int8_w[41] = (|vec_data_041_d2);
    mask_d2_int8_w[42] = (|vec_data_042_d2);
    mask_d2_int8_w[43] = (|vec_data_043_d2);
    mask_d2_int8_w[44] = (|vec_data_044_d2);
    mask_d2_int8_w[45] = (|vec_data_045_d2);
    mask_d2_int8_w[46] = (|vec_data_046_d2);
    mask_d2_int8_w[47] = (|vec_data_047_d2);
    mask_d2_int8_w[48] = (|vec_data_048_d2);
    mask_d2_int8_w[49] = (|vec_data_049_d2);
    mask_d2_int8_w[50] = (|vec_data_050_d2);
    mask_d2_int8_w[51] = (|vec_data_051_d2);
    mask_d2_int8_w[52] = (|vec_data_052_d2);
    mask_d2_int8_w[53] = (|vec_data_053_d2);
    mask_d2_int8_w[54] = (|vec_data_054_d2);
    mask_d2_int8_w[55] = (|vec_data_055_d2);
    mask_d2_int8_w[56] = (|vec_data_056_d2);
    mask_d2_int8_w[57] = (|vec_data_057_d2);
    mask_d2_int8_w[58] = (|vec_data_058_d2);
    mask_d2_int8_w[59] = (|vec_data_059_d2);
    mask_d2_int8_w[60] = (|vec_data_060_d2);
    mask_d2_int8_w[61] = (|vec_data_061_d2);
    mask_d2_int8_w[62] = (|vec_data_062_d2);
    mask_d2_int8_w[63] = (|vec_data_063_d2);
    mask_d2_int8_w[64] = (|vec_data_064_d2);
    mask_d2_int8_w[65] = (|vec_data_065_d2);
    mask_d2_int8_w[66] = (|vec_data_066_d2);
    mask_d2_int8_w[67] = (|vec_data_067_d2);
    mask_d2_int8_w[68] = (|vec_data_068_d2);
    mask_d2_int8_w[69] = (|vec_data_069_d2);
    mask_d2_int8_w[70] = (|vec_data_070_d2);
    mask_d2_int8_w[71] = (|vec_data_071_d2);
    mask_d2_int8_w[72] = (|vec_data_072_d2);
    mask_d2_int8_w[73] = (|vec_data_073_d2);
    mask_d2_int8_w[74] = (|vec_data_074_d2);
    mask_d2_int8_w[75] = (|vec_data_075_d2);
    mask_d2_int8_w[76] = (|vec_data_076_d2);
    mask_d2_int8_w[77] = (|vec_data_077_d2);
    mask_d2_int8_w[78] = (|vec_data_078_d2);
    mask_d2_int8_w[79] = (|vec_data_079_d2);
    mask_d2_int8_w[80] = (|vec_data_080_d2);
    mask_d2_int8_w[81] = (|vec_data_081_d2);
    mask_d2_int8_w[82] = (|vec_data_082_d2);
    mask_d2_int8_w[83] = (|vec_data_083_d2);
    mask_d2_int8_w[84] = (|vec_data_084_d2);
    mask_d2_int8_w[85] = (|vec_data_085_d2);
    mask_d2_int8_w[86] = (|vec_data_086_d2);
    mask_d2_int8_w[87] = (|vec_data_087_d2);
    mask_d2_int8_w[88] = (|vec_data_088_d2);
    mask_d2_int8_w[89] = (|vec_data_089_d2);
    mask_d2_int8_w[90] = (|vec_data_090_d2);
    mask_d2_int8_w[91] = (|vec_data_091_d2);
    mask_d2_int8_w[92] = (|vec_data_092_d2);
    mask_d2_int8_w[93] = (|vec_data_093_d2);
    mask_d2_int8_w[94] = (|vec_data_094_d2);
    mask_d2_int8_w[95] = (|vec_data_095_d2);
    mask_d2_int8_w[96] = (|vec_data_096_d2);
    mask_d2_int8_w[97] = (|vec_data_097_d2);
    mask_d2_int8_w[98] = (|vec_data_098_d2);
    mask_d2_int8_w[99] = (|vec_data_099_d2);
    mask_d2_int8_w[100] = (|vec_data_100_d2);
    mask_d2_int8_w[101] = (|vec_data_101_d2);
    mask_d2_int8_w[102] = (|vec_data_102_d2);
    mask_d2_int8_w[103] = (|vec_data_103_d2);
    mask_d2_int8_w[104] = (|vec_data_104_d2);
    mask_d2_int8_w[105] = (|vec_data_105_d2);
    mask_d2_int8_w[106] = (|vec_data_106_d2);
    mask_d2_int8_w[107] = (|vec_data_107_d2);
    mask_d2_int8_w[108] = (|vec_data_108_d2);
    mask_d2_int8_w[109] = (|vec_data_109_d2);
    mask_d2_int8_w[110] = (|vec_data_110_d2);
    mask_d2_int8_w[111] = (|vec_data_111_d2);
    mask_d2_int8_w[112] = (|vec_data_112_d2);
    mask_d2_int8_w[113] = (|vec_data_113_d2);
    mask_d2_int8_w[114] = (|vec_data_114_d2);
    mask_d2_int8_w[115] = (|vec_data_115_d2);
    mask_d2_int8_w[116] = (|vec_data_116_d2);
    mask_d2_int8_w[117] = (|vec_data_117_d2);
    mask_d2_int8_w[118] = (|vec_data_118_d2);
    mask_d2_int8_w[119] = (|vec_data_119_d2);
    mask_d2_int8_w[120] = (|vec_data_120_d2);
    mask_d2_int8_w[121] = (|vec_data_121_d2);
    mask_d2_int8_w[122] = (|vec_data_122_d2);
    mask_d2_int8_w[123] = (|vec_data_123_d2);
    mask_d2_int8_w[124] = (|vec_data_124_d2);
    mask_d2_int8_w[125] = (|vec_data_125_d2);
    mask_d2_int8_w[126] = (|vec_data_126_d2);
    mask_d2_int8_w[127] = (|vec_data_127_d2);
end


always @(
  vec_data_001_d2
  or vec_data_000_d2
  or vec_data_003_d2
  or vec_data_002_d2
  or vec_data_005_d2
  or vec_data_004_d2
  or vec_data_007_d2
  or vec_data_006_d2
  or vec_data_009_d2
  or vec_data_008_d2
  or vec_data_011_d2
  or vec_data_010_d2
  or vec_data_013_d2
  or vec_data_012_d2
  or vec_data_015_d2
  or vec_data_014_d2
  or vec_data_017_d2
  or vec_data_016_d2
  or vec_data_019_d2
  or vec_data_018_d2
  or vec_data_021_d2
  or vec_data_020_d2
  or vec_data_023_d2
  or vec_data_022_d2
  or vec_data_025_d2
  or vec_data_024_d2
  or vec_data_027_d2
  or vec_data_026_d2
  or vec_data_029_d2
  or vec_data_028_d2
  or vec_data_031_d2
  or vec_data_030_d2
  or vec_data_033_d2
  or vec_data_032_d2
  or vec_data_035_d2
  or vec_data_034_d2
  or vec_data_037_d2
  or vec_data_036_d2
  or vec_data_039_d2
  or vec_data_038_d2
  or vec_data_041_d2
  or vec_data_040_d2
  or vec_data_043_d2
  or vec_data_042_d2
  or vec_data_045_d2
  or vec_data_044_d2
  or vec_data_047_d2
  or vec_data_046_d2
  or vec_data_049_d2
  or vec_data_048_d2
  or vec_data_051_d2
  or vec_data_050_d2
  or vec_data_053_d2
  or vec_data_052_d2
  or vec_data_055_d2
  or vec_data_054_d2
  or vec_data_057_d2
  or vec_data_056_d2
  or vec_data_059_d2
  or vec_data_058_d2
  or vec_data_061_d2
  or vec_data_060_d2
  or vec_data_063_d2
  or vec_data_062_d2
  or vec_data_065_d2
  or vec_data_064_d2
  or vec_data_067_d2
  or vec_data_066_d2
  or vec_data_069_d2
  or vec_data_068_d2
  or vec_data_071_d2
  or vec_data_070_d2
  or vec_data_073_d2
  or vec_data_072_d2
  or vec_data_075_d2
  or vec_data_074_d2
  or vec_data_077_d2
  or vec_data_076_d2
  or vec_data_079_d2
  or vec_data_078_d2
  or vec_data_081_d2
  or vec_data_080_d2
  or vec_data_083_d2
  or vec_data_082_d2
  or vec_data_085_d2
  or vec_data_084_d2
  or vec_data_087_d2
  or vec_data_086_d2
  or vec_data_089_d2
  or vec_data_088_d2
  or vec_data_091_d2
  or vec_data_090_d2
  or vec_data_093_d2
  or vec_data_092_d2
  or vec_data_095_d2
  or vec_data_094_d2
  or vec_data_097_d2
  or vec_data_096_d2
  or vec_data_099_d2
  or vec_data_098_d2
  or vec_data_101_d2
  or vec_data_100_d2
  or vec_data_103_d2
  or vec_data_102_d2
  or vec_data_105_d2
  or vec_data_104_d2
  or vec_data_107_d2
  or vec_data_106_d2
  or vec_data_109_d2
  or vec_data_108_d2
  or vec_data_111_d2
  or vec_data_110_d2
  or vec_data_113_d2
  or vec_data_112_d2
  or vec_data_115_d2
  or vec_data_114_d2
  or vec_data_117_d2
  or vec_data_116_d2
  or vec_data_119_d2
  or vec_data_118_d2
  or vec_data_121_d2
  or vec_data_120_d2
  or vec_data_123_d2
  or vec_data_122_d2
  or vec_data_125_d2
  or vec_data_124_d2
  or vec_data_127_d2
  or vec_data_126_d2
  ) begin
    mask_d2_int16_w[1:0] = {2{(|{vec_data_001_d2, vec_data_000_d2})}};
    mask_d2_int16_w[3:2] = {2{(|{vec_data_003_d2, vec_data_002_d2})}};
    mask_d2_int16_w[5:4] = {2{(|{vec_data_005_d2, vec_data_004_d2})}};
    mask_d2_int16_w[7:6] = {2{(|{vec_data_007_d2, vec_data_006_d2})}};
    mask_d2_int16_w[9:8] = {2{(|{vec_data_009_d2, vec_data_008_d2})}};
    mask_d2_int16_w[11:10] = {2{(|{vec_data_011_d2, vec_data_010_d2})}};
    mask_d2_int16_w[13:12] = {2{(|{vec_data_013_d2, vec_data_012_d2})}};
    mask_d2_int16_w[15:14] = {2{(|{vec_data_015_d2, vec_data_014_d2})}};
    mask_d2_int16_w[17:16] = {2{(|{vec_data_017_d2, vec_data_016_d2})}};
    mask_d2_int16_w[19:18] = {2{(|{vec_data_019_d2, vec_data_018_d2})}};
    mask_d2_int16_w[21:20] = {2{(|{vec_data_021_d2, vec_data_020_d2})}};
    mask_d2_int16_w[23:22] = {2{(|{vec_data_023_d2, vec_data_022_d2})}};
    mask_d2_int16_w[25:24] = {2{(|{vec_data_025_d2, vec_data_024_d2})}};
    mask_d2_int16_w[27:26] = {2{(|{vec_data_027_d2, vec_data_026_d2})}};
    mask_d2_int16_w[29:28] = {2{(|{vec_data_029_d2, vec_data_028_d2})}};
    mask_d2_int16_w[31:30] = {2{(|{vec_data_031_d2, vec_data_030_d2})}};
    mask_d2_int16_w[33:32] = {2{(|{vec_data_033_d2, vec_data_032_d2})}};
    mask_d2_int16_w[35:34] = {2{(|{vec_data_035_d2, vec_data_034_d2})}};
    mask_d2_int16_w[37:36] = {2{(|{vec_data_037_d2, vec_data_036_d2})}};
    mask_d2_int16_w[39:38] = {2{(|{vec_data_039_d2, vec_data_038_d2})}};
    mask_d2_int16_w[41:40] = {2{(|{vec_data_041_d2, vec_data_040_d2})}};
    mask_d2_int16_w[43:42] = {2{(|{vec_data_043_d2, vec_data_042_d2})}};
    mask_d2_int16_w[45:44] = {2{(|{vec_data_045_d2, vec_data_044_d2})}};
    mask_d2_int16_w[47:46] = {2{(|{vec_data_047_d2, vec_data_046_d2})}};
    mask_d2_int16_w[49:48] = {2{(|{vec_data_049_d2, vec_data_048_d2})}};
    mask_d2_int16_w[51:50] = {2{(|{vec_data_051_d2, vec_data_050_d2})}};
    mask_d2_int16_w[53:52] = {2{(|{vec_data_053_d2, vec_data_052_d2})}};
    mask_d2_int16_w[55:54] = {2{(|{vec_data_055_d2, vec_data_054_d2})}};
    mask_d2_int16_w[57:56] = {2{(|{vec_data_057_d2, vec_data_056_d2})}};
    mask_d2_int16_w[59:58] = {2{(|{vec_data_059_d2, vec_data_058_d2})}};
    mask_d2_int16_w[61:60] = {2{(|{vec_data_061_d2, vec_data_060_d2})}};
    mask_d2_int16_w[63:62] = {2{(|{vec_data_063_d2, vec_data_062_d2})}};
    mask_d2_int16_w[65:64] = {2{(|{vec_data_065_d2, vec_data_064_d2})}};
    mask_d2_int16_w[67:66] = {2{(|{vec_data_067_d2, vec_data_066_d2})}};
    mask_d2_int16_w[69:68] = {2{(|{vec_data_069_d2, vec_data_068_d2})}};
    mask_d2_int16_w[71:70] = {2{(|{vec_data_071_d2, vec_data_070_d2})}};
    mask_d2_int16_w[73:72] = {2{(|{vec_data_073_d2, vec_data_072_d2})}};
    mask_d2_int16_w[75:74] = {2{(|{vec_data_075_d2, vec_data_074_d2})}};
    mask_d2_int16_w[77:76] = {2{(|{vec_data_077_d2, vec_data_076_d2})}};
    mask_d2_int16_w[79:78] = {2{(|{vec_data_079_d2, vec_data_078_d2})}};
    mask_d2_int16_w[81:80] = {2{(|{vec_data_081_d2, vec_data_080_d2})}};
    mask_d2_int16_w[83:82] = {2{(|{vec_data_083_d2, vec_data_082_d2})}};
    mask_d2_int16_w[85:84] = {2{(|{vec_data_085_d2, vec_data_084_d2})}};
    mask_d2_int16_w[87:86] = {2{(|{vec_data_087_d2, vec_data_086_d2})}};
    mask_d2_int16_w[89:88] = {2{(|{vec_data_089_d2, vec_data_088_d2})}};
    mask_d2_int16_w[91:90] = {2{(|{vec_data_091_d2, vec_data_090_d2})}};
    mask_d2_int16_w[93:92] = {2{(|{vec_data_093_d2, vec_data_092_d2})}};
    mask_d2_int16_w[95:94] = {2{(|{vec_data_095_d2, vec_data_094_d2})}};
    mask_d2_int16_w[97:96] = {2{(|{vec_data_097_d2, vec_data_096_d2})}};
    mask_d2_int16_w[99:98] = {2{(|{vec_data_099_d2, vec_data_098_d2})}};
    mask_d2_int16_w[101:100] = {2{(|{vec_data_101_d2, vec_data_100_d2})}};
    mask_d2_int16_w[103:102] = {2{(|{vec_data_103_d2, vec_data_102_d2})}};
    mask_d2_int16_w[105:104] = {2{(|{vec_data_105_d2, vec_data_104_d2})}};
    mask_d2_int16_w[107:106] = {2{(|{vec_data_107_d2, vec_data_106_d2})}};
    mask_d2_int16_w[109:108] = {2{(|{vec_data_109_d2, vec_data_108_d2})}};
    mask_d2_int16_w[111:110] = {2{(|{vec_data_111_d2, vec_data_110_d2})}};
    mask_d2_int16_w[113:112] = {2{(|{vec_data_113_d2, vec_data_112_d2})}};
    mask_d2_int16_w[115:114] = {2{(|{vec_data_115_d2, vec_data_114_d2})}};
    mask_d2_int16_w[117:116] = {2{(|{vec_data_117_d2, vec_data_116_d2})}};
    mask_d2_int16_w[119:118] = {2{(|{vec_data_119_d2, vec_data_118_d2})}};
    mask_d2_int16_w[121:120] = {2{(|{vec_data_121_d2, vec_data_120_d2})}};
    mask_d2_int16_w[123:122] = {2{(|{vec_data_123_d2, vec_data_122_d2})}};
    mask_d2_int16_w[125:124] = {2{(|{vec_data_125_d2, vec_data_124_d2})}};
    mask_d2_int16_w[127:126] = {2{(|{vec_data_127_d2, vec_data_126_d2})}};
end


always @(
  vec_data_001_d2
  or vec_data_000_d2
  or vec_data_003_d2
  or vec_data_002_d2
  or vec_data_005_d2
  or vec_data_004_d2
  or vec_data_007_d2
  or vec_data_006_d2
  or vec_data_009_d2
  or vec_data_008_d2
  or vec_data_011_d2
  or vec_data_010_d2
  or vec_data_013_d2
  or vec_data_012_d2
  or vec_data_015_d2
  or vec_data_014_d2
  or vec_data_017_d2
  or vec_data_016_d2
  or vec_data_019_d2
  or vec_data_018_d2
  or vec_data_021_d2
  or vec_data_020_d2
  or vec_data_023_d2
  or vec_data_022_d2
  or vec_data_025_d2
  or vec_data_024_d2
  or vec_data_027_d2
  or vec_data_026_d2
  or vec_data_029_d2
  or vec_data_028_d2
  or vec_data_031_d2
  or vec_data_030_d2
  or vec_data_033_d2
  or vec_data_032_d2
  or vec_data_035_d2
  or vec_data_034_d2
  or vec_data_037_d2
  or vec_data_036_d2
  or vec_data_039_d2
  or vec_data_038_d2
  or vec_data_041_d2
  or vec_data_040_d2
  or vec_data_043_d2
  or vec_data_042_d2
  or vec_data_045_d2
  or vec_data_044_d2
  or vec_data_047_d2
  or vec_data_046_d2
  or vec_data_049_d2
  or vec_data_048_d2
  or vec_data_051_d2
  or vec_data_050_d2
  or vec_data_053_d2
  or vec_data_052_d2
  or vec_data_055_d2
  or vec_data_054_d2
  or vec_data_057_d2
  or vec_data_056_d2
  or vec_data_059_d2
  or vec_data_058_d2
  or vec_data_061_d2
  or vec_data_060_d2
  or vec_data_063_d2
  or vec_data_062_d2
  or vec_data_065_d2
  or vec_data_064_d2
  or vec_data_067_d2
  or vec_data_066_d2
  or vec_data_069_d2
  or vec_data_068_d2
  or vec_data_071_d2
  or vec_data_070_d2
  or vec_data_073_d2
  or vec_data_072_d2
  or vec_data_075_d2
  or vec_data_074_d2
  or vec_data_077_d2
  or vec_data_076_d2
  or vec_data_079_d2
  or vec_data_078_d2
  or vec_data_081_d2
  or vec_data_080_d2
  or vec_data_083_d2
  or vec_data_082_d2
  or vec_data_085_d2
  or vec_data_084_d2
  or vec_data_087_d2
  or vec_data_086_d2
  or vec_data_089_d2
  or vec_data_088_d2
  or vec_data_091_d2
  or vec_data_090_d2
  or vec_data_093_d2
  or vec_data_092_d2
  or vec_data_095_d2
  or vec_data_094_d2
  or vec_data_097_d2
  or vec_data_096_d2
  or vec_data_099_d2
  or vec_data_098_d2
  or vec_data_101_d2
  or vec_data_100_d2
  or vec_data_103_d2
  or vec_data_102_d2
  or vec_data_105_d2
  or vec_data_104_d2
  or vec_data_107_d2
  or vec_data_106_d2
  or vec_data_109_d2
  or vec_data_108_d2
  or vec_data_111_d2
  or vec_data_110_d2
  or vec_data_113_d2
  or vec_data_112_d2
  or vec_data_115_d2
  or vec_data_114_d2
  or vec_data_117_d2
  or vec_data_116_d2
  or vec_data_119_d2
  or vec_data_118_d2
  or vec_data_121_d2
  or vec_data_120_d2
  or vec_data_123_d2
  or vec_data_122_d2
  or vec_data_125_d2
  or vec_data_124_d2
  or vec_data_127_d2
  or vec_data_126_d2
  ) begin
    mask_d2_fp16_w[1:0] = {2{(|{vec_data_001_d2[6:0], vec_data_000_d2})}};
    mask_d2_fp16_w[3:2] = {2{(|{vec_data_003_d2[6:0], vec_data_002_d2})}};
    mask_d2_fp16_w[5:4] = {2{(|{vec_data_005_d2[6:0], vec_data_004_d2})}};
    mask_d2_fp16_w[7:6] = {2{(|{vec_data_007_d2[6:0], vec_data_006_d2})}};
    mask_d2_fp16_w[9:8] = {2{(|{vec_data_009_d2[6:0], vec_data_008_d2})}};
    mask_d2_fp16_w[11:10] = {2{(|{vec_data_011_d2[6:0], vec_data_010_d2})}};
    mask_d2_fp16_w[13:12] = {2{(|{vec_data_013_d2[6:0], vec_data_012_d2})}};
    mask_d2_fp16_w[15:14] = {2{(|{vec_data_015_d2[6:0], vec_data_014_d2})}};
    mask_d2_fp16_w[17:16] = {2{(|{vec_data_017_d2[6:0], vec_data_016_d2})}};
    mask_d2_fp16_w[19:18] = {2{(|{vec_data_019_d2[6:0], vec_data_018_d2})}};
    mask_d2_fp16_w[21:20] = {2{(|{vec_data_021_d2[6:0], vec_data_020_d2})}};
    mask_d2_fp16_w[23:22] = {2{(|{vec_data_023_d2[6:0], vec_data_022_d2})}};
    mask_d2_fp16_w[25:24] = {2{(|{vec_data_025_d2[6:0], vec_data_024_d2})}};
    mask_d2_fp16_w[27:26] = {2{(|{vec_data_027_d2[6:0], vec_data_026_d2})}};
    mask_d2_fp16_w[29:28] = {2{(|{vec_data_029_d2[6:0], vec_data_028_d2})}};
    mask_d2_fp16_w[31:30] = {2{(|{vec_data_031_d2[6:0], vec_data_030_d2})}};
    mask_d2_fp16_w[33:32] = {2{(|{vec_data_033_d2[6:0], vec_data_032_d2})}};
    mask_d2_fp16_w[35:34] = {2{(|{vec_data_035_d2[6:0], vec_data_034_d2})}};
    mask_d2_fp16_w[37:36] = {2{(|{vec_data_037_d2[6:0], vec_data_036_d2})}};
    mask_d2_fp16_w[39:38] = {2{(|{vec_data_039_d2[6:0], vec_data_038_d2})}};
    mask_d2_fp16_w[41:40] = {2{(|{vec_data_041_d2[6:0], vec_data_040_d2})}};
    mask_d2_fp16_w[43:42] = {2{(|{vec_data_043_d2[6:0], vec_data_042_d2})}};
    mask_d2_fp16_w[45:44] = {2{(|{vec_data_045_d2[6:0], vec_data_044_d2})}};
    mask_d2_fp16_w[47:46] = {2{(|{vec_data_047_d2[6:0], vec_data_046_d2})}};
    mask_d2_fp16_w[49:48] = {2{(|{vec_data_049_d2[6:0], vec_data_048_d2})}};
    mask_d2_fp16_w[51:50] = {2{(|{vec_data_051_d2[6:0], vec_data_050_d2})}};
    mask_d2_fp16_w[53:52] = {2{(|{vec_data_053_d2[6:0], vec_data_052_d2})}};
    mask_d2_fp16_w[55:54] = {2{(|{vec_data_055_d2[6:0], vec_data_054_d2})}};
    mask_d2_fp16_w[57:56] = {2{(|{vec_data_057_d2[6:0], vec_data_056_d2})}};
    mask_d2_fp16_w[59:58] = {2{(|{vec_data_059_d2[6:0], vec_data_058_d2})}};
    mask_d2_fp16_w[61:60] = {2{(|{vec_data_061_d2[6:0], vec_data_060_d2})}};
    mask_d2_fp16_w[63:62] = {2{(|{vec_data_063_d2[6:0], vec_data_062_d2})}};
    mask_d2_fp16_w[65:64] = {2{(|{vec_data_065_d2[6:0], vec_data_064_d2})}};
    mask_d2_fp16_w[67:66] = {2{(|{vec_data_067_d2[6:0], vec_data_066_d2})}};
    mask_d2_fp16_w[69:68] = {2{(|{vec_data_069_d2[6:0], vec_data_068_d2})}};
    mask_d2_fp16_w[71:70] = {2{(|{vec_data_071_d2[6:0], vec_data_070_d2})}};
    mask_d2_fp16_w[73:72] = {2{(|{vec_data_073_d2[6:0], vec_data_072_d2})}};
    mask_d2_fp16_w[75:74] = {2{(|{vec_data_075_d2[6:0], vec_data_074_d2})}};
    mask_d2_fp16_w[77:76] = {2{(|{vec_data_077_d2[6:0], vec_data_076_d2})}};
    mask_d2_fp16_w[79:78] = {2{(|{vec_data_079_d2[6:0], vec_data_078_d2})}};
    mask_d2_fp16_w[81:80] = {2{(|{vec_data_081_d2[6:0], vec_data_080_d2})}};
    mask_d2_fp16_w[83:82] = {2{(|{vec_data_083_d2[6:0], vec_data_082_d2})}};
    mask_d2_fp16_w[85:84] = {2{(|{vec_data_085_d2[6:0], vec_data_084_d2})}};
    mask_d2_fp16_w[87:86] = {2{(|{vec_data_087_d2[6:0], vec_data_086_d2})}};
    mask_d2_fp16_w[89:88] = {2{(|{vec_data_089_d2[6:0], vec_data_088_d2})}};
    mask_d2_fp16_w[91:90] = {2{(|{vec_data_091_d2[6:0], vec_data_090_d2})}};
    mask_d2_fp16_w[93:92] = {2{(|{vec_data_093_d2[6:0], vec_data_092_d2})}};
    mask_d2_fp16_w[95:94] = {2{(|{vec_data_095_d2[6:0], vec_data_094_d2})}};
    mask_d2_fp16_w[97:96] = {2{(|{vec_data_097_d2[6:0], vec_data_096_d2})}};
    mask_d2_fp16_w[99:98] = {2{(|{vec_data_099_d2[6:0], vec_data_098_d2})}};
    mask_d2_fp16_w[101:100] = {2{(|{vec_data_101_d2[6:0], vec_data_100_d2})}};
    mask_d2_fp16_w[103:102] = {2{(|{vec_data_103_d2[6:0], vec_data_102_d2})}};
    mask_d2_fp16_w[105:104] = {2{(|{vec_data_105_d2[6:0], vec_data_104_d2})}};
    mask_d2_fp16_w[107:106] = {2{(|{vec_data_107_d2[6:0], vec_data_106_d2})}};
    mask_d2_fp16_w[109:108] = {2{(|{vec_data_109_d2[6:0], vec_data_108_d2})}};
    mask_d2_fp16_w[111:110] = {2{(|{vec_data_111_d2[6:0], vec_data_110_d2})}};
    mask_d2_fp16_w[113:112] = {2{(|{vec_data_113_d2[6:0], vec_data_112_d2})}};
    mask_d2_fp16_w[115:114] = {2{(|{vec_data_115_d2[6:0], vec_data_114_d2})}};
    mask_d2_fp16_w[117:116] = {2{(|{vec_data_117_d2[6:0], vec_data_116_d2})}};
    mask_d2_fp16_w[119:118] = {2{(|{vec_data_119_d2[6:0], vec_data_118_d2})}};
    mask_d2_fp16_w[121:120] = {2{(|{vec_data_121_d2[6:0], vec_data_120_d2})}};
    mask_d2_fp16_w[123:122] = {2{(|{vec_data_123_d2[6:0], vec_data_122_d2})}};
    mask_d2_fp16_w[125:124] = {2{(|{vec_data_125_d2[6:0], vec_data_124_d2})}};
    mask_d2_fp16_w[127:126] = {2{(|{vec_data_127_d2[6:0], vec_data_126_d2})}};
end


always @(
  is_int8
  or mask_d2_int8_w
  or is_fp16
  or mask_d2_fp16_w
  or mask_d2_int16_w
  ) begin
    mask_d2_w = is_int8 ? mask_d2_int8_w :
                is_fp16 ? mask_d2_fp16_w :
                mask_d2_int16_w;
end


always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    valid_d3 <= 1'b0;
  end else begin
  valid_d3 <= valid_d2;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    mask_d3 <= mask_d2_w;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    mask_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    sel_d3 <= sel_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    sel_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_000_d3 <= vec_data_000_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_000_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_001_d3 <= vec_data_001_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_001_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_002_d3 <= vec_data_002_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_002_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_003_d3 <= vec_data_003_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_003_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_004_d3 <= vec_data_004_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_004_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_005_d3 <= vec_data_005_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_005_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_006_d3 <= vec_data_006_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_006_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_007_d3 <= vec_data_007_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_007_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_008_d3 <= vec_data_008_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_008_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_009_d3 <= vec_data_009_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_009_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_010_d3 <= vec_data_010_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_010_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_011_d3 <= vec_data_011_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_011_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_012_d3 <= vec_data_012_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_012_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_013_d3 <= vec_data_013_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_013_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_014_d3 <= vec_data_014_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_014_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_015_d3 <= vec_data_015_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_015_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_016_d3 <= vec_data_016_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_016_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_017_d3 <= vec_data_017_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_017_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_018_d3 <= vec_data_018_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_018_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_019_d3 <= vec_data_019_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_019_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_020_d3 <= vec_data_020_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_020_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_021_d3 <= vec_data_021_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_021_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_022_d3 <= vec_data_022_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_022_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_023_d3 <= vec_data_023_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_023_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_024_d3 <= vec_data_024_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_024_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_025_d3 <= vec_data_025_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_025_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_026_d3 <= vec_data_026_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_026_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_027_d3 <= vec_data_027_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_027_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_028_d3 <= vec_data_028_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_028_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_029_d3 <= vec_data_029_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_029_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_030_d3 <= vec_data_030_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_030_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_031_d3 <= vec_data_031_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_031_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_032_d3 <= vec_data_032_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_032_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_033_d3 <= vec_data_033_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_033_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_034_d3 <= vec_data_034_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_034_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_035_d3 <= vec_data_035_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_035_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_036_d3 <= vec_data_036_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_036_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_037_d3 <= vec_data_037_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_037_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_038_d3 <= vec_data_038_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_038_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_039_d3 <= vec_data_039_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_039_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_040_d3 <= vec_data_040_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_040_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_041_d3 <= vec_data_041_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_041_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_042_d3 <= vec_data_042_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_042_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_043_d3 <= vec_data_043_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_043_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_044_d3 <= vec_data_044_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_044_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_045_d3 <= vec_data_045_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_045_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_046_d3 <= vec_data_046_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_046_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_047_d3 <= vec_data_047_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_047_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_048_d3 <= vec_data_048_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_048_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_049_d3 <= vec_data_049_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_049_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_050_d3 <= vec_data_050_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_050_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_051_d3 <= vec_data_051_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_051_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_052_d3 <= vec_data_052_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_052_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_053_d3 <= vec_data_053_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_053_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_054_d3 <= vec_data_054_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_054_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_055_d3 <= vec_data_055_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_055_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_056_d3 <= vec_data_056_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_056_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_057_d3 <= vec_data_057_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_057_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_058_d3 <= vec_data_058_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_058_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_059_d3 <= vec_data_059_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_059_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_060_d3 <= vec_data_060_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_060_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_061_d3 <= vec_data_061_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_061_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_062_d3 <= vec_data_062_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_062_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_063_d3 <= vec_data_063_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_063_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_064_d3 <= vec_data_064_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_064_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_065_d3 <= vec_data_065_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_065_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_066_d3 <= vec_data_066_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_066_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_067_d3 <= vec_data_067_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_067_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_068_d3 <= vec_data_068_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_068_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_069_d3 <= vec_data_069_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_069_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_070_d3 <= vec_data_070_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_070_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_071_d3 <= vec_data_071_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_071_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_072_d3 <= vec_data_072_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_072_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_073_d3 <= vec_data_073_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_073_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_074_d3 <= vec_data_074_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_074_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_075_d3 <= vec_data_075_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_075_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_076_d3 <= vec_data_076_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_076_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_077_d3 <= vec_data_077_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_077_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_078_d3 <= vec_data_078_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_078_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_079_d3 <= vec_data_079_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_079_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_080_d3 <= vec_data_080_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_080_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_081_d3 <= vec_data_081_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_081_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_082_d3 <= vec_data_082_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_082_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_083_d3 <= vec_data_083_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_083_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_084_d3 <= vec_data_084_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_084_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_085_d3 <= vec_data_085_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_085_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_086_d3 <= vec_data_086_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_086_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_087_d3 <= vec_data_087_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_087_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_088_d3 <= vec_data_088_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_088_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_089_d3 <= vec_data_089_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_089_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_090_d3 <= vec_data_090_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_090_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_091_d3 <= vec_data_091_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_091_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_092_d3 <= vec_data_092_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_092_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_093_d3 <= vec_data_093_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_093_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_094_d3 <= vec_data_094_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_094_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_095_d3 <= vec_data_095_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_095_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_096_d3 <= vec_data_096_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_096_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_097_d3 <= vec_data_097_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_097_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_098_d3 <= vec_data_098_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_098_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_099_d3 <= vec_data_099_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_099_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_100_d3 <= vec_data_100_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_100_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_101_d3 <= vec_data_101_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_101_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_102_d3 <= vec_data_102_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_102_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_103_d3 <= vec_data_103_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_103_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_104_d3 <= vec_data_104_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_104_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_105_d3 <= vec_data_105_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_105_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_106_d3 <= vec_data_106_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_106_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_107_d3 <= vec_data_107_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_107_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_108_d3 <= vec_data_108_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_108_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_109_d3 <= vec_data_109_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_109_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_110_d3 <= vec_data_110_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_110_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_111_d3 <= vec_data_111_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_111_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_112_d3 <= vec_data_112_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_112_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_113_d3 <= vec_data_113_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_113_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_114_d3 <= vec_data_114_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_114_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_115_d3 <= vec_data_115_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_115_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_116_d3 <= vec_data_116_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_116_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_117_d3 <= vec_data_117_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_117_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_118_d3 <= vec_data_118_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_118_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_119_d3 <= vec_data_119_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_119_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_120_d3 <= vec_data_120_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_120_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_121_d3 <= vec_data_121_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_121_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_122_d3 <= vec_data_122_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_122_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_123_d3 <= vec_data_123_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_123_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_124_d3 <= vec_data_124_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_124_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_125_d3 <= vec_data_125_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_125_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_126_d3 <= vec_data_126_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_126_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((valid_d2) == 1'b1) begin
    vec_data_127_d3 <= vec_data_127_d2;
  // VCS coverage off
  end else if ((valid_d2) == 1'b0) begin
  end else begin
    vec_data_127_d3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


////////////////////////////////// output: rename //////////////////////////////////
assign output_pvld = valid_d3;
assign output_mask = mask_d3;
assign output_sel = sel_d3;
assign output_data0 = vec_data_000_d3;
assign output_data1 = vec_data_001_d3;
assign output_data2 = vec_data_002_d3;
assign output_data3 = vec_data_003_d3;
assign output_data4 = vec_data_004_d3;
assign output_data5 = vec_data_005_d3;
assign output_data6 = vec_data_006_d3;
assign output_data7 = vec_data_007_d3;
assign output_data8 = vec_data_008_d3;
assign output_data9 = vec_data_009_d3;
assign output_data10 = vec_data_010_d3;
assign output_data11 = vec_data_011_d3;
assign output_data12 = vec_data_012_d3;
assign output_data13 = vec_data_013_d3;
assign output_data14 = vec_data_014_d3;
assign output_data15 = vec_data_015_d3;
assign output_data16 = vec_data_016_d3;
assign output_data17 = vec_data_017_d3;
assign output_data18 = vec_data_018_d3;
assign output_data19 = vec_data_019_d3;
assign output_data20 = vec_data_020_d3;
assign output_data21 = vec_data_021_d3;
assign output_data22 = vec_data_022_d3;
assign output_data23 = vec_data_023_d3;
assign output_data24 = vec_data_024_d3;
assign output_data25 = vec_data_025_d3;
assign output_data26 = vec_data_026_d3;
assign output_data27 = vec_data_027_d3;
assign output_data28 = vec_data_028_d3;
assign output_data29 = vec_data_029_d3;
assign output_data30 = vec_data_030_d3;
assign output_data31 = vec_data_031_d3;
assign output_data32 = vec_data_032_d3;
assign output_data33 = vec_data_033_d3;
assign output_data34 = vec_data_034_d3;
assign output_data35 = vec_data_035_d3;
assign output_data36 = vec_data_036_d3;
assign output_data37 = vec_data_037_d3;
assign output_data38 = vec_data_038_d3;
assign output_data39 = vec_data_039_d3;
assign output_data40 = vec_data_040_d3;
assign output_data41 = vec_data_041_d3;
assign output_data42 = vec_data_042_d3;
assign output_data43 = vec_data_043_d3;
assign output_data44 = vec_data_044_d3;
assign output_data45 = vec_data_045_d3;
assign output_data46 = vec_data_046_d3;
assign output_data47 = vec_data_047_d3;
assign output_data48 = vec_data_048_d3;
assign output_data49 = vec_data_049_d3;
assign output_data50 = vec_data_050_d3;
assign output_data51 = vec_data_051_d3;
assign output_data52 = vec_data_052_d3;
assign output_data53 = vec_data_053_d3;
assign output_data54 = vec_data_054_d3;
assign output_data55 = vec_data_055_d3;
assign output_data56 = vec_data_056_d3;
assign output_data57 = vec_data_057_d3;
assign output_data58 = vec_data_058_d3;
assign output_data59 = vec_data_059_d3;
assign output_data60 = vec_data_060_d3;
assign output_data61 = vec_data_061_d3;
assign output_data62 = vec_data_062_d3;
assign output_data63 = vec_data_063_d3;
assign output_data64 = vec_data_064_d3;
assign output_data65 = vec_data_065_d3;
assign output_data66 = vec_data_066_d3;
assign output_data67 = vec_data_067_d3;
assign output_data68 = vec_data_068_d3;
assign output_data69 = vec_data_069_d3;
assign output_data70 = vec_data_070_d3;
assign output_data71 = vec_data_071_d3;
assign output_data72 = vec_data_072_d3;
assign output_data73 = vec_data_073_d3;
assign output_data74 = vec_data_074_d3;
assign output_data75 = vec_data_075_d3;
assign output_data76 = vec_data_076_d3;
assign output_data77 = vec_data_077_d3;
assign output_data78 = vec_data_078_d3;
assign output_data79 = vec_data_079_d3;
assign output_data80 = vec_data_080_d3;
assign output_data81 = vec_data_081_d3;
assign output_data82 = vec_data_082_d3;
assign output_data83 = vec_data_083_d3;
assign output_data84 = vec_data_084_d3;
assign output_data85 = vec_data_085_d3;
assign output_data86 = vec_data_086_d3;
assign output_data87 = vec_data_087_d3;
assign output_data88 = vec_data_088_d3;
assign output_data89 = vec_data_089_d3;
assign output_data90 = vec_data_090_d3;
assign output_data91 = vec_data_091_d3;
assign output_data92 = vec_data_092_d3;
assign output_data93 = vec_data_093_d3;
assign output_data94 = vec_data_094_d3;
assign output_data95 = vec_data_095_d3;
assign output_data96 = vec_data_096_d3;
assign output_data97 = vec_data_097_d3;
assign output_data98 = vec_data_098_d3;
assign output_data99 = vec_data_099_d3;
assign output_data100 = vec_data_100_d3;
assign output_data101 = vec_data_101_d3;
assign output_data102 = vec_data_102_d3;
assign output_data103 = vec_data_103_d3;
assign output_data104 = vec_data_104_d3;
assign output_data105 = vec_data_105_d3;
assign output_data106 = vec_data_106_d3;
assign output_data107 = vec_data_107_d3;
assign output_data108 = vec_data_108_d3;
assign output_data109 = vec_data_109_d3;
assign output_data110 = vec_data_110_d3;
assign output_data111 = vec_data_111_d3;
assign output_data112 = vec_data_112_d3;
assign output_data113 = vec_data_113_d3;
assign output_data114 = vec_data_114_d3;
assign output_data115 = vec_data_115_d3;
assign output_data116 = vec_data_116_d3;
assign output_data117 = vec_data_117_d3;
assign output_data118 = vec_data_118_d3;
assign output_data119 = vec_data_119_d3;
assign output_data120 = vec_data_120_d3;
assign output_data121 = vec_data_121_d3;
assign output_data122 = vec_data_122_d3;
assign output_data123 = vec_data_123_d3;
assign output_data124 = vec_data_124_d3;
assign output_data125 = vec_data_125_d3;
assign output_data126 = vec_data_126_d3;
assign output_data127 = vec_data_127_d3;



endmodule // NV_NVDLA_CSC_WL_dec


