`ifndef _MEM_DEFINE_SVH
`define _MEM_DEFINE_SVH

  `define MEM_ADDR_WIDTH    32

`endif
