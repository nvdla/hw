`ifndef _CSB_DEFINES_SVH_
`define _CSB_DEFINES_SVH_

//-------------------------------------------------------------------------------------
//
// MACROS: csb defines
//
// XXX
//-------------------------------------------------------------------------------------

`ifndef CSB_ADDR_WIDTH
`define CSB_ADDR_WIDTH 16
`endif

`ifndef CSB_DATA_WIDTH
`define CSB_DATA_WIDTH 32
`endif

`endif // _CSB_DEFINES_SVH_
