//
// Component: XXX
//
// Description:
/// @file 
/// XXX
//

module nvdla_tg_top;
    
    initial begin
      	run_test("nvdla_tg_base_test");
    end

endmodule
