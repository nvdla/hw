// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

//nvdla_top sv side SC-SV Adapter 
// This is autogenerated code */

`ifndef _nvdla_top_sv_layer
`define _nvdla_top_sv_layer

//////////////////////////////////////////////////////
// Callback Header file
//////////////////////////////////////////////////////
//Include nvdla_top_sv_tlm_callbacks.svh 
//for callback classes. They are declared, constructed and registered
// via the nvdla_top_DEC_MACRO, nvdla_top_CONSTRUCT_MACRO and nvdla_top_REGISTER_MACRO
// defined in nvdla_top_sv_tlm_callbacks.svh
`ifdef nvdla_top_NEED_SCSV_SV_CALLBACKS
`include "nvdla_top_sv_tlm_callbacks.svh"
`endif

class nvdla_top_sv_layer extends uvm_component;

    `uvm_component_utils(nvdla_top_sv_layer)

    /////////////////////////////////////////////////////////
    //TLM Connector Proxy and Passthrough Socket Declaration
    /////////////////////////////////////////////////////////
 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt; //initiator passthrough for nvdla_core2dbb_axi4 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sc2sv_nvdla_core2dbb_axi4; //Connector Proxy for nvdla_core2dbb_axi4 
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt; //initiator passthrough for nvdla_core2cvsram_axi4 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sc2sv_nvdla_core2cvsram_axi4; //Connector Proxy for nvdla_core2cvsram_axi4 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sc2sv_dma_monitor_cv; //Connector Proxy for dma_monitor_cv
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_dma_monitor_cv_initiator_pt; //initiator passthrough for dma_monitor_cv
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sv2sc_dma_monitor_cv_credit; //Connector Proxy for dma_monitor_cv_credit
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt; //target passthrough for dma_monitor_cv_credit
`endif
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_nvdla_host_master_if_target_pt; //target passthrough for nvdla_host_master_if 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sv2sc_nvdla_host_master_if; //Connector Proxy for nvdla_host_master_if 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_dma_monitor_mc_initiator_pt; //initiator passthrough for dma_monitor_mc 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sc2sv_dma_monitor_mc; //Connector Proxy for dma_monitor_mc 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt; //initiator passthrough for convolution_core_monitor_initiator 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sc2sv_convolution_core_monitor_initiator; //Connector Proxy for convolution_core_monitor_initiator 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt; //initiator passthrough for post_processing_monitor_initiator 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sc2sv_post_processing_monitor_initiator; //Connector Proxy for post_processing_monitor_initiator 
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt; //target passthrough for dma_monitor_mc_credit 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sv2sc_dma_monitor_mc_credit; //Connector Proxy for dma_monitor_mc_credit 
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt; //target passthrough for convolution_core_monitor_credit 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sv2sc_convolution_core_monitor_credit; //Connector Proxy for convolution_core_monitor_credit 
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_post_processing_monitor_credit_target_pt; //target passthrough for post_processing_monitor_credit 
    nvdla_scsv_sv_tlm_channel #(tlm_generic_payload) nvdla_top_sv2sc_post_processing_monitor_credit; //Connector Proxy for post_processing_monitor_credit  

    //nvdla_top Virtual Interface
    virtual nvdla_top_sv_interface nvdla_top_sv_interface_inst;

    ///////////////////////////////////////////////////////////////////////////
    //Callback declaration
    //This macro expands to the declaration lines of the callback classes
    //This is expected to be defined in nvdla_top_sv_tlm_callbacks.svh
`ifdef nvdla_top_DEC_MACRO
    `nvdla_top_DEC_MACRO

`endif

    /////////////////////////////////////////////////////////////
    //// constructor
    /////////////////////////////////////////////////////////////
    function new(string name, uvm_component parent = null);
        super.new(name, parent);
    endfunction // new
    
      
    /////////////////////////////////////////////////////////////
    /// build phase()
    /////////////////////////////////////////////////////////////
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        /////////////////////////////////////////////////////////
        //TLM Connector Proxy and Passthrough Socket Construction
        /////////////////////////////////////////////////////////     
        nvdla_top_sc2sv_nvdla_core2dbb_axi4 = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_nvdla_core2dbb_axi4",this); 
        nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt = new ("nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt",this);     
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
        nvdla_top_sc2sv_nvdla_core2cvsram_axi4 = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_nvdla_core2cvsram_axi4",this); 
        nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt = new ("nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt",this);     
        nvdla_top_sc2sv_dma_monitor_cv = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_dma_monitor_cv",this);
        nvdla_top_sc2sv_dma_monitor_cv_initiator_pt = new ("nvdla_top_sc2sv_dma_monitor_cv_initiator_pt",this);
        nvdla_top_sv2sc_dma_monitor_cv_credit = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_dma_monitor_cv_credit",this);
        nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt = new ("nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt",this);
`endif
        nvdla_top_sv2sc_nvdla_host_master_if = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_nvdla_host_master_if",this); 
        nvdla_top_sv2sc_nvdla_host_master_if_target_pt = new ("nvdla_top_sv2sc_nvdla_host_master_if_target_pt",this);     
        nvdla_top_sc2sv_dma_monitor_mc = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_dma_monitor_mc",this); 
        nvdla_top_sc2sv_dma_monitor_mc_initiator_pt = new ("nvdla_top_sc2sv_dma_monitor_mc_initiator_pt",this);     
        nvdla_top_sc2sv_convolution_core_monitor_initiator = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_convolution_core_monitor_initiator",this); 
        nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt = new ("nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt",this);     
        nvdla_top_sc2sv_post_processing_monitor_initiator = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sc2sv_post_processing_monitor_initiator",this); 
        nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt = new ("nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt",this);     
        nvdla_top_sv2sc_dma_monitor_mc_credit = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_dma_monitor_mc_credit",this); 
        nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt = new ("nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt",this);     
        nvdla_top_sv2sc_convolution_core_monitor_credit = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_convolution_core_monitor_credit",this); 
        nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt = new ("nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt",this);     
        nvdla_top_sv2sc_post_processing_monitor_credit = nvdla_scsv_sv_tlm_channel#(tlm_generic_payload)::type_id::create("nvdla_top_sv2sc_post_processing_monitor_credit",this); 
        nvdla_top_sv2sc_post_processing_monitor_credit_target_pt = new ("nvdla_top_sv2sc_post_processing_monitor_credit_target_pt",this);  

        ///////////////////////////////////////////////////////////////////////////
        //Callback Construction
        //This macro expands to the construction calls for the callback classes
        //This is expected to be defined in nvdla_top_sv_tlm_callbacks.svh
`ifdef nvdla_top_CONSTRUCT_MACRO
        `nvdla_top_CONSTRUCT_MACRO

`endif

    endfunction : build_phase
    
      
    /////////////////////////////////////////////////////////////
    /// connect phase()
    /////////////////////////////////////////////////////////////
    virtual function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);

             
        /////////////////////////////////////////////////////////////
        /// Get nvdla_top interface handle from uvm_config_db
        /////////////////////////////////////////////////////////////
        if (!uvm_config_db#(virtual nvdla_top_sv_interface)::get(this, "", "nvdla_top_sv_interface", nvdla_top_sv_interface_inst)) begin
            `uvm_fatal({get_name(),"/NO_VIF"},"No Interface found to connect signals to");
        end

        ////////////////////////////////////////////////////////////////////////////////////////////
        /// Hierarchial TLM connections from connector proxies to respective passthrough sockets
        ////////////////////////////////////////////////////////////////////////////////////////////

        nvdla_top_sc2sv_nvdla_core2dbb_axi4.sv_tlm_initiator.connect(nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sc2sv_nvdla_core2dbb_axi4.sv_tlm_target, "nvdla_top_sc2sv_nvdla_core2dbb_axi4");
         
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
        nvdla_top_sc2sv_nvdla_core2cvsram_axi4.sv_tlm_initiator.connect(nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sc2sv_nvdla_core2cvsram_axi4.sv_tlm_target, "nvdla_top_sc2sv_nvdla_core2cvsram_axi4");
        nvdla_top_sc2sv_dma_monitor_cv.sv_tlm_initiator.connect(nvdla_top_sc2sv_dma_monitor_cv_initiator_pt);
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sc2sv_dma_monitor_cv.sv_tlm_target, "nvdla_top_sc2sv_dma_monitor_cv");
        nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt.connect(nvdla_top_sv2sc_dma_monitor_cv_credit.sv_tlm_target);
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sv2sc_dma_monitor_cv_credit.sv_tlm_initiator, "nvdla_top_sv2sc_dma_monitor_cv_credit");
`endif
         
        nvdla_top_sv2sc_nvdla_host_master_if_target_pt.connect(nvdla_top_sv2sc_nvdla_host_master_if.sv_tlm_target);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sv2sc_nvdla_host_master_if.sv_tlm_initiator, "nvdla_top_sv2sc_nvdla_host_master_if"); 
        nvdla_top_sc2sv_dma_monitor_mc.sv_tlm_initiator.connect(nvdla_top_sc2sv_dma_monitor_mc_initiator_pt);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sc2sv_dma_monitor_mc.sv_tlm_target, "nvdla_top_sc2sv_dma_monitor_mc");
         
         
        nvdla_top_sc2sv_convolution_core_monitor_initiator.sv_tlm_initiator.connect(nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sc2sv_convolution_core_monitor_initiator.sv_tlm_target, "nvdla_top_sc2sv_convolution_core_monitor_initiator");
         
        nvdla_top_sc2sv_post_processing_monitor_initiator.sv_tlm_initiator.connect(nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sc2sv_post_processing_monitor_initiator.sv_tlm_target, "nvdla_top_sc2sv_post_processing_monitor_initiator");
         
        nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt.connect(nvdla_top_sv2sc_dma_monitor_mc_credit.sv_tlm_target);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sv2sc_dma_monitor_mc_credit.sv_tlm_initiator, "nvdla_top_sv2sc_dma_monitor_mc_credit"); 
        nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt.connect(nvdla_top_sv2sc_convolution_core_monitor_credit.sv_tlm_target);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sv2sc_convolution_core_monitor_credit.sv_tlm_initiator, "nvdla_top_sv2sc_convolution_core_monitor_credit"); 
        nvdla_top_sv2sc_post_processing_monitor_credit_target_pt.connect(nvdla_top_sv2sc_post_processing_monitor_credit.sv_tlm_target);               
        uvmc_tlm #(.T(tlm_generic_payload),.CVRT(nvdla_scsv_converter))::connect(nvdla_top_sv2sc_post_processing_monitor_credit.sv_tlm_initiator, "nvdla_top_sv2sc_post_processing_monitor_credit"); 

        ///////////////////////////////////////////////////////////////////////////
        //Callback Registration
        //This macro expands to the registration calls(::add) for the callback classes
        //This is expected to be defined in nvdla_top_sv_tlm_callbacks.svh
`ifdef nvdla_top_REGISTER_MACRO
        `nvdla_top_REGISTER_MACRO

`endif 
    endfunction : connect_phase

endclass:nvdla_top_sv_layer

`endif // nvdla_top_sv_layer 
