`ifndef _DP_DEFINES_SV_
`define _DP_DEFINES_SV_



`endif // _DP_DEFINES_SV_
