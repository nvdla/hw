// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_NVDLA_RT_cacc2glb.v

module NV_NVDLA_RT_cacc2glb (
   nvdla_core_clk
  ,nvdla_core_rstn
  ,cacc2glb_done_intr_src_pd
  ,cacc2glb_done_intr_dst_pd
  );

//
// NV_NVDLA_RT_cacc2glb_ports.v
// DO NOT EDIT, generated by ness version 2.0, backend=verilog
//
// Command: /home/ip/shared/inf/ness/2.0/38823533/bin/run_ispec_backend verilog nvdla_all.nessdb defs.touch-verilog -backend_opt '--nogenerate_io_capture' -backend_opt '--generate_ports'
input  nvdla_core_clk;
input  nvdla_core_rstn;

//<-- cacc2glb_done_intr_src clk=nvdla_core_clk flow=none ctype=nvdla_glb_intr_source_t c_hdr=nvdla_glb_intr_source_iface.h
input [1:0] cacc2glb_done_intr_src_pd;

output [1:0] cacc2glb_done_intr_dst_pd;

wire [1:0] cacc2glb_done_intr_pd_d0;
reg  [1:0] cacc2glb_done_intr_pd_d1;
reg  [1:0] cacc2glb_done_intr_pd_d2;



assign cacc2glb_done_intr_pd_d0 = cacc2glb_done_intr_src_pd;


always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    cacc2glb_done_intr_pd_d1 <= {2{1'b0}};
  end else begin
  cacc2glb_done_intr_pd_d1 <= cacc2glb_done_intr_pd_d0;
  end
end


always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    cacc2glb_done_intr_pd_d2 <= {2{1'b0}};
  end else begin
  cacc2glb_done_intr_pd_d2 <= cacc2glb_done_intr_pd_d1;
  end
end


assign cacc2glb_done_intr_dst_pd = cacc2glb_done_intr_pd_d2;



endmodule // NV_NVDLA_RT_cacc2glb

