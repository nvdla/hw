`ifndef _NVDLA_TG_BASE_TEST_SV_
`define _NVDLA_TG_BASE_TEST_SV_

//-------------------------------------------------------------------------------------
//
// CLASS: nvdla_tg_base_test 
//
// @description: this is the test base of all user defined trace generator tests
//-------------------------------------------------------------------------------------

`include "nvdla_tg_core.sv"
class nvdla_tg_base_test extends uvm_test;

    string                      inst_name;
    /*
        layers: number of layers to be generated by current test
    */
    int                         layers;
     /*
        cur_test_layer: counter of how many times generator is active, e.g. gets called by test
    */
    int                         cur_test_layer;
   
    int                         fh;
    /*
        generator: trace generator instance
    */
    nvdla_tg_core               generator;  
    
    /*
        Methods
    */
    extern function new(string name="nvdla_base_test", uvm_component parent);
    extern function set_inst_name(string inst_name=""); 
    /*
        override_scenario_pool: handle for user defined test to manipulate scenario pool.
        by default no override is enabled
        if per-layer override is required, please use along with variable cur_test_layer
    */
    extern virtual function override_scenario_pool();
    extern         function void pre_abort();
    extern         function void do_report();
    /*
        Phases
    */
    extern function void end_of_elaboration_phase(uvm_phase phase);
    extern task          main_phase(uvm_phase phase);
    extern function void report_phase(uvm_phase phase);
    
    `uvm_component_utils_begin(nvdla_tg_base_test)
        `uvm_field_int(layers, UVM_ALL_ON)
    `uvm_component_utils_end

endclass : nvdla_tg_base_test

function nvdla_tg_base_test::new(string name="nvdla_base_test", uvm_component parent);
    super.new(name,parent);
    generator = nvdla_tg_core::type_id::create("TRACE_GENERATOR", this);
    fh = 0;
    layers = 1;
endfunction:new

function nvdla_tg_base_test::set_inst_name(string inst_name="");
    this.inst_name = inst_name;
endfunction: set_inst_name

function void nvdla_tg_base_test::end_of_elaboration_phase(uvm_phase phase);
    super.end_of_elaboration_phase(phase);

    begin
        uvm_factory factory = uvm_factory::get();
        factory.print();
        uvm_top.print_topology();
    end
endfunction: end_of_elaboration_phase

task nvdla_tg_base_test::main_phase(uvm_phase phase);
    `uvm_info(inst_name, $sformatf("main_phase begins ..."), UVM_HIGH)
    phase.raise_objection(this);
    
    fh = $fopen({inst_name.tolower(),".cfg"});
    if(fh==0) begin
        `uvm_fatal(inst_name,"Fail to create trace file ...");
    end else begin
        `uvm_info(inst_name,$sformatf("Create trace file %s ...",{inst_name.tolower(),"_autogen_trace"}),UVM_LOW);
    end
    
    if(layers==0) begin
        `uvm_fatal(inst_name, "Please explictly specify a layer number via command line ...");
    end

    for(cur_test_layer=0;cur_test_layer<layers;cur_test_layer++) begin
        generator.restore_scenario_pool();
        override_scenario_pool();
        generator.generate_trace(fh);
    end
    $fclose(fh);

    `uvm_info(inst_name, $sformatf("main_phase finishes ..."), UVM_HIGH)
    phase.drop_objection(this);
endtask: main_phase

function nvdla_tg_base_test::override_scenario_pool();
    `uvm_info(inst_name, "No scenario override ...", UVM_HIGH);
endfunction: override_scenario_pool

function void nvdla_tg_base_test::report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info(inst_name, $sformatf("report_phase begin ..."), UVM_HIGH)

    do_report();
endfunction : report_phase

function void nvdla_tg_base_test::pre_abort();
    super.pre_abort();
    do_report();
endfunction

// Added for post-processing
function void nvdla_tg_base_test::do_report();
    uvm_report_server rs = uvm_report_server::get_server();
    if (rs.get_severity_count(UVM_FATAL) + rs.get_severity_count(UVM_ERROR) == 0) begin
        $display("*****************************");
        $display("**  TRACE GENERATION PASS  **");
        $display("*****************************");
    end else begin
        $display("*****************************");
        $display("**  TRACE GENERATION FAIL  **");
        $display("*****************************");
    end
endfunction

`endif //_NVDLA_TG_BASE_TEST_SV_
