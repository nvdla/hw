
// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: nvdla_top_config.tt






//This is autogenerated code
//This is the layer component
//IP Name nvdla_top
//Filename nvdla_top_sv_adapter

`ifndef _nvdla_top_sv_adapter
`define _nvdla_top_sv_adapter

class nvdla_top_sv_adapter extends uvm_component;

    `uvm_component_utils(nvdla_top_sv_adapter)
    /////////////////////////////////////////////////////////////
    // Passthrough TLM sockets declaration
    /////////////////////////////////////////////////////////////
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt; 
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt; 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_dma_monitor_cv_initiator_pt;
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt;
`endif
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_nvdla_host_master_if_target_pt; 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_dma_monitor_mc_initiator_pt; 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt; 
    uvm_tlm_b_passthrough_initiator_socket#(tlm_generic_payload) nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt; 
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt; 
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt; 
    uvm_tlm_b_passthrough_target_socket#(tlm_generic_payload) nvdla_top_sv2sc_post_processing_monitor_credit_target_pt;  


    /////////////////////////////////////////////////////////////
    // Layer component instantiation
    /////////////////////////////////////////////////////////////
    nvdla_top_sv_layer nvdla_top_sv_layer_inst;

    /////////////////////////////////////////////////////////////
    //// constructor
    /////////////////////////////////////////////////////////////
    function new(string name, uvm_component parent = null);
        super.new(name, parent);
    endfunction // new
    
      
    /////////////////////////////////////////////////////////////
    /// build phase()
    /////////////////////////////////////////////////////////////
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        /////////////////////////////////////////////////////////
        //Layer Construction
         ///////////////////////////////////////////////////////// 
        nvdla_top_sv_layer_inst = nvdla_top_sv_layer::type_id::create("nvdla_top_sv_layer_inst",this);

        /////////////////////////////////////////////////////////
        //Passthrough Socket Construction
        ///////////////////////////////////////////////////////// 
         nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt = new ("nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt",this); 
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
         nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt = new ("nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt",this); 
         nvdla_top_sc2sv_dma_monitor_cv_initiator_pt = new ("nvdla_top_sc2sv_dma_monitor_cv_initiator_pt",this);
         nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt = new ("nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt",this);
`endif
         nvdla_top_sv2sc_nvdla_host_master_if_target_pt = new ("nvdla_top_sv2sc_nvdla_host_master_if_target_pt",this); 
         nvdla_top_sc2sv_dma_monitor_mc_initiator_pt = new ("nvdla_top_sc2sv_dma_monitor_mc_initiator_pt",this); 
         nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt = new ("nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt",this); 
         nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt = new ("nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt",this); 
         nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt = new ("nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt",this); 
         nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt = new ("nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt",this); 
         nvdla_top_sv2sc_post_processing_monitor_credit_target_pt = new ("nvdla_top_sv2sc_post_processing_monitor_credit_target_pt",this);  
        //////////////////////////////////////////////////////////////////////
        //  Instantiate user converters
        //////////////////////////////////////////////////////////////////////


    endfunction : build_phase
    
      
    /////////////////////////////////////////////////////////////
    /// connect phase()
    /////////////////////////////////////////////////////////////
    virtual function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);

        ////////////////////////////////////////////////////////////////////////////////////////////
        // Connect sockets to SC side via UVM-Connect calls
        // Hierarchial TLM connection from layer's passthrough sockets to adapter passthrough sockets 
        ////////////////////////////////////////////////////////////////////////////////////////////
         nvdla_top_sv_layer_inst.nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt.connect(nvdla_top_sc2sv_nvdla_core2dbb_axi4_initiator_pt);
         
`ifdef NVDLA_SECONDARY_MEMIF_ENABLE
         nvdla_top_sv_layer_inst.nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt.connect(nvdla_top_sc2sv_nvdla_core2cvsram_axi4_initiator_pt);
         nvdla_top_sv_layer_inst.nvdla_top_sc2sv_dma_monitor_cv_initiator_pt.connect(nvdla_top_sc2sv_dma_monitor_cv_initiator_pt);
         nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt.connect(nvdla_top_sv_layer_inst.nvdla_top_sv2sc_dma_monitor_cv_credit_target_pt);
`endif         
         nvdla_top_sv2sc_nvdla_host_master_if_target_pt.connect(nvdla_top_sv_layer_inst.nvdla_top_sv2sc_nvdla_host_master_if_target_pt);
         nvdla_top_sv_layer_inst.nvdla_top_sc2sv_dma_monitor_mc_initiator_pt.connect(nvdla_top_sc2sv_dma_monitor_mc_initiator_pt);
         
         
         nvdla_top_sv_layer_inst.nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt.connect(nvdla_top_sc2sv_convolution_core_monitor_initiator_initiator_pt);
         
         nvdla_top_sv_layer_inst.nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt.connect(nvdla_top_sc2sv_post_processing_monitor_initiator_initiator_pt);
         
         nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt.connect(nvdla_top_sv_layer_inst.nvdla_top_sv2sc_dma_monitor_mc_credit_target_pt);
         nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt.connect(nvdla_top_sv_layer_inst.nvdla_top_sv2sc_convolution_core_monitor_credit_target_pt);
         nvdla_top_sv2sc_post_processing_monitor_credit_target_pt.connect(nvdla_top_sv_layer_inst.nvdla_top_sv2sc_post_processing_monitor_credit_target_pt); 

    endfunction : connect_phase


endclass:nvdla_top_sv_adapter

`endif // nvdla_top_sv_adapter 
