// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_NVDLA_SDP_CORE_Y_core.v

module SDP_Y_CORE_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_CORE_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module SDP_Y_CORE_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_CORE_mgc_io_sync_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module SDP_Y_CORE_mgc_io_sync_v1 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


module SDP_Y_CORE_mgc_in_sync_v1 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v4.v 
module SDP_Y_CORE_mgc_shift_bl_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SIGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ../td_ccore_solutions/leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-136
//  Generated date: Fri Jun 16 21:48:25 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_leading_sign_49_0
// ------------------------------------------------------------------


module SDP_Y_CORE_leading_sign_49_0 (
  mantissa, rtn
);
  input [48:0] mantissa;
  output [5:0] rtn;


  // Interconnect Declarations
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_22;
  wire c_h_1_23;

  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[42:41]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[34:33]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = (mantissa[26:25]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = (mantissa[18:17]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 & c_h_1_12 & c_h_1_13;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = (mantissa[10:9]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = (mantissa[2:1]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (c_h_1_22
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = c_h_1_6 & (c_h_1_13 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4)) & (~((~(c_h_1_21
      & (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4))) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = c_h_1_2 & (c_h_1_5 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3)) & (~((~(c_h_1_9
      & (c_h_1_12 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~(((~(c_h_1_17 & (c_h_1_20 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2)) & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~(((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2)))) & c_h_1_21))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl
      = ((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01))))) & (~(((mantissa[44])
      | (~((mantissa[43:42]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))))
      & (~(((mantissa[36]) | (~((mantissa[35:34]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01))))) & (~(((mantissa[28])
      | (~((mantissa[27:26]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))))
      & (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~(((~((~((mantissa[16]) | (~((mantissa[15:14]!=2'b01))))) &
      (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[8])
      | (~((mantissa[7:6]!=2'b01))))) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)))) | c_h_1_22) & c_h_1_23))) | ((~ (mantissa[0]))
      & c_h_1_22 & c_h_1_23);
  assign rtn = {c_h_1_23 , (IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl)};
endmodule




//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v 
module SDP_Y_CORE_mgc_shift_l_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_CORE_mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module SDP_Y_CORE_mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v4.v 
module SDP_Y_CORE_mgc_shift_r_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_out_fifo_wait_core_v2001_v9.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module SDP_Y_CORE_mgc_out_fifo_wait_core_v9 (clk, en, arst, srst, ld, vd, d, lz, vz,  z, sd);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer ph_clk  =  1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en   =  1; // clock enable polarity
    parameter integer ph_arst =  1; // async reset polarity
    parameter integer ph_srst =  1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)

   localparam integer  fifo_b = width * fifo_sz;

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;
    output    [sz_width-1:0]      sd; 

    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;
    reg      [fifo_mx:0] stat_pre;
    reg      [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    wire     [fifo_mx:0] en_l;
    wire     [fifo_mx_over_8:0] en_l_s;

    reg       [width-1:0] buff_nxt;

    reg                   stat_nxt;
    reg                   stat_before;
    reg                   stat_after;
    reg       [fifo_mx:0] en_l_var;

    integer               i;
    genvar                eni;

    wire [32:0]           size_t;
    reg [31:0]            count;
    reg [31:0]            count_t;
    reg [32:0]            n_elem;
    // synopsys translate_off
    reg [31:0]            peak = 32'b0;
    // synopsys translate_on
    wire                  active;

    assign active = ld | vz; // (ld & ~vd) | (vz & ~lz);

    genvar igen;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      wire [31:0]           delta;
      //  0 :  32'b0      if ld==0 and (vz & stat[fifo_sz-1])==0   
      //               or if ld==1 and (vz & stat[fifo_sz-1])==1
      // +1 :  32'b1      if ld==1 and (vz & stat[fifo_sz-1])==0
      // -1 : {32{1'b1}}  if ld==0 and (vz & stat[fifo_sz-1])==1
      assign delta   =  {{31{(~ld & (vz & stat[fifo_sz-1]))}} , (vz & stat[fifo_sz-1]) ^ ld};
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = count + delta;
      assign sd = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_before = (i != 0) ? stat[i-1] : 1'b0;
          stat_after = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;
          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));
  
          stat_pre[i] = stat_nxt;
          if (vz & stat_before )
            begin
              buff_nxt[0+:width] = buff[width*(i-1)+:width];
              en_l_var[i] = 1'b1;
            end
          else if (ld & ~((~vz) & stat[i]))
            begin
              buff_nxt = d;
              en_l_var[i] = 1'b1;
            end
          else
            begin
              buff_nxt = d; // Don't care input to disabled flop
              en_l_var[i] = 1'b0;
            end
             
          buff_pre[width*i+:width] = buff_nxt[0+:width];
  
          if ((stat_after == 1'b1) & (stat[i] == 1'b0)) 
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end

        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else 
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        if ( peak < count )
          peak = count;
        // synopsys translate_on
      end

      if (ph_en) begin: PH_EN_HI
        assign en_l_s[fifo_mx_over_8] = en & active;
        for (igen = 0 ; igen < fifo_sz ; igen = igen + 1) begin: NEED_A_LABEL
          assign en_l[igen] = en & en_l_var[igen];
        end
        for (igen = 1 ; igen <= fifo_mx_over_8 ; igen = igen + 1) begin: NEED_A_LABEL2
          assign  en_l_s[igen-1] = en & (stat[igen*8]) & (active);
        end
      end
      else begin: PH_EN_LO
        assign en_l_s[fifo_mx_over_8] = en | ~active;
        for (igen = 0 ; igen < fifo_sz ; igen = igen + 1) begin: NEED_A_LABEL3
          assign en_l[igen] = en | ~en_l_var[igen];
        end
        for (igen = 1 ; igen <= fifo_mx_over_8 ; igen = igen + 1) begin: NEED_A_LABEL2
          assign  en_l_s[igen-1] = en | (~stat[igen*8]) | (~active);
        end
      end

      // Output registers:
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: BUF_GEN
        if (ph_clk==1) begin: POS_BUF
          if (ph_arst==0) begin: LABEL1
            always @(posedge clk or negedge arst)
            if (arst == 1'b0) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
          else begin: LABEL2 // ph_arst==1
            always @(posedge clk or posedge arst)
            if (arst == 1'b1) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
        end
        else begin: NEG_BUF
          if (ph_arst==0) begin: LABEL3
            always @(negedge clk or negedge arst)
            if (arst == 1'b0) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
          else begin: LABEL4 // ph_arst==1
            always @(negedge clk or posedge arst)
            if (arst == 1'b1) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
        end
      end

      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: STATGEN2
        if (ph_clk==1) begin: POS_STAT
          if (ph_arst==0) begin: LABEL5
            always @(posedge clk or negedge arst)
            if (arst == 1'b0) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
          else begin: LABEL6 // ph_arst==1
            always @(posedge clk or posedge arst)
            if (arst == 1'b1) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
        end
        else begin: NEG_STAT // ph_clk==0
          if (ph_arst==0) begin: LABEL7
            always @(negedge clk or negedge arst)
            if (arst == 1'b0) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
          else begin: LABEL8 // ph_arst==1
            always @(negedge clk or posedge arst)
            if (arst == 1'b1) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign sd = ld & ~vz;
    end
    endgenerate

endmodule



//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_pipe_v2001_v10.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 *
 *    vdout - can be considered as a notFULL signal
 *    vdin  - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from ldout & !vdout
 *    read_stall  - an internal debug signal formed from ldin & !vdin
 *
 */
// two clock pipe
module SDP_Y_CORE_mgc_pipe_v10 (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, sd);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter integer ph_clk  = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en   = 1;  // clock enable polarity
    parameter integer ph_arst = 1;  // async reset polarity
    parameter integer ph_srst = 1;  // sync reset polarity

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output [sz_width-1:0]      sd;

    // synopsys translate_off
    wire               write_stall;
    wire               read_stall;
    assign write_stall = ldout & !vdout;
    assign read_stall = ldin & !vdin;
    // synopsys translate_on

    SDP_Y_CORE_mgc_out_fifo_wait_core_v9
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (vdin),
        .vz      (ldin),
        .z       (din),
        .sd      (sd)
    );

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-159
//  Generated date: Mon Jul  3 19:09:52 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_truncate_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_truncate_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_mul_op_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_mul_op_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_mul_src_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_mul_src_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_mul_prelu_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_mul_prelu_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_mul_bypass_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_mul_bypass_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_chn_mul_out_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_chn_mul_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_chn_mul_op_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_chn_mul_op_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_chn_mul_in_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_chn_mul_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for Y_mul_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : Y_mul_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_staller
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_mul_in_rsci_wen_comp, core_wten,
      chn_mul_op_rsci_wen_comp, chn_mul_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_mul_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_mul_op_rsci_wen_comp;
  input chn_mul_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_mul_in_rsci_wen_comp & chn_mul_op_rsci_wen_comp & chn_mul_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_truncate_rsc_triosy_obj_bawt, cfg_truncate_rsc_triosy_obj_biwt,
      cfg_truncate_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_truncate_rsc_triosy_obj_bawt;
  input cfg_truncate_rsc_triosy_obj_biwt;
  input cfg_truncate_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_truncate_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_truncate_rsc_triosy_obj_bawt = cfg_truncate_rsc_triosy_obj_biwt | cfg_truncate_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_truncate_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_truncate_rsc_triosy_obj_bcwt <= ~((~(cfg_truncate_rsc_triosy_obj_bcwt |
          cfg_truncate_rsc_triosy_obj_biwt)) | cfg_truncate_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_ctrl (
  cfg_truncate_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_truncate_rsc_triosy_obj_iswt0,
      cfg_truncate_rsc_triosy_obj_biwt, cfg_truncate_rsc_triosy_obj_bdwt
);
  input cfg_truncate_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_truncate_rsc_triosy_obj_iswt0;
  output cfg_truncate_rsc_triosy_obj_biwt;
  output cfg_truncate_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_truncate_rsc_triosy_obj_biwt = (~ core_wten) & cfg_truncate_rsc_triosy_obj_iswt0;
  assign cfg_truncate_rsc_triosy_obj_bdwt = cfg_truncate_rsc_triosy_obj_oswt & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_op_rsc_triosy_obj_bawt, cfg_mul_op_rsc_triosy_obj_biwt,
      cfg_mul_op_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_op_rsc_triosy_obj_bawt;
  input cfg_mul_op_rsc_triosy_obj_biwt;
  input cfg_mul_op_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_mul_op_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_op_rsc_triosy_obj_bawt = cfg_mul_op_rsc_triosy_obj_biwt | cfg_mul_op_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_op_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_op_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_op_rsc_triosy_obj_bcwt | cfg_mul_op_rsc_triosy_obj_biwt))
          | cfg_mul_op_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl (
  cfg_mul_op_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_op_rsc_triosy_obj_iswt0,
      cfg_mul_op_rsc_triosy_obj_biwt, cfg_mul_op_rsc_triosy_obj_bdwt
);
  input cfg_mul_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_op_rsc_triosy_obj_iswt0;
  output cfg_mul_op_rsc_triosy_obj_biwt;
  output cfg_mul_op_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_op_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_op_rsc_triosy_obj_iswt0;
  assign cfg_mul_op_rsc_triosy_obj_bdwt = cfg_mul_op_rsc_triosy_obj_oswt & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_src_rsc_triosy_obj_bawt, cfg_mul_src_rsc_triosy_obj_biwt,
      cfg_mul_src_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_src_rsc_triosy_obj_bawt;
  input cfg_mul_src_rsc_triosy_obj_biwt;
  input cfg_mul_src_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_mul_src_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_src_rsc_triosy_obj_bawt = cfg_mul_src_rsc_triosy_obj_biwt | cfg_mul_src_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_src_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_src_rsc_triosy_obj_bcwt | cfg_mul_src_rsc_triosy_obj_biwt))
          | cfg_mul_src_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl (
  cfg_mul_src_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_src_rsc_triosy_obj_iswt0,
      cfg_mul_src_rsc_triosy_obj_biwt, cfg_mul_src_rsc_triosy_obj_bdwt
);
  input cfg_mul_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_src_rsc_triosy_obj_iswt0;
  output cfg_mul_src_rsc_triosy_obj_biwt;
  output cfg_mul_src_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_src_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_src_rsc_triosy_obj_iswt0;
  assign cfg_mul_src_rsc_triosy_obj_bdwt = cfg_mul_src_rsc_triosy_obj_oswt & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_prelu_rsc_triosy_obj_bawt, cfg_mul_prelu_rsc_triosy_obj_biwt,
      cfg_mul_prelu_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_prelu_rsc_triosy_obj_bawt;
  input cfg_mul_prelu_rsc_triosy_obj_biwt;
  input cfg_mul_prelu_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_mul_prelu_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_prelu_rsc_triosy_obj_bawt = cfg_mul_prelu_rsc_triosy_obj_biwt |
      cfg_mul_prelu_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_prelu_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_prelu_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_prelu_rsc_triosy_obj_bcwt
          | cfg_mul_prelu_rsc_triosy_obj_biwt)) | cfg_mul_prelu_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl
    (
  cfg_mul_prelu_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_prelu_rsc_triosy_obj_iswt0,
      cfg_mul_prelu_rsc_triosy_obj_biwt, cfg_mul_prelu_rsc_triosy_obj_bdwt
);
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_prelu_rsc_triosy_obj_iswt0;
  output cfg_mul_prelu_rsc_triosy_obj_biwt;
  output cfg_mul_prelu_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_prelu_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_prelu_rsc_triosy_obj_iswt0;
  assign cfg_mul_prelu_rsc_triosy_obj_bdwt = cfg_mul_prelu_rsc_triosy_obj_oswt &
      core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_bypass_rsc_triosy_obj_bawt, cfg_mul_bypass_rsc_triosy_obj_biwt,
      cfg_mul_bypass_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_bypass_rsc_triosy_obj_bawt;
  input cfg_mul_bypass_rsc_triosy_obj_biwt;
  input cfg_mul_bypass_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_mul_bypass_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_bypass_rsc_triosy_obj_bawt = cfg_mul_bypass_rsc_triosy_obj_biwt
      | cfg_mul_bypass_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_bypass_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_mul_bypass_rsc_triosy_obj_bcwt <= ~((~(cfg_mul_bypass_rsc_triosy_obj_bcwt
          | cfg_mul_bypass_rsc_triosy_obj_biwt)) | cfg_mul_bypass_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl
    (
  cfg_mul_bypass_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_mul_bypass_rsc_triosy_obj_iswt0,
      cfg_mul_bypass_rsc_triosy_obj_biwt, cfg_mul_bypass_rsc_triosy_obj_bdwt
);
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_bypass_rsc_triosy_obj_iswt0;
  output cfg_mul_bypass_rsc_triosy_obj_biwt;
  output cfg_mul_bypass_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_mul_bypass_rsc_triosy_obj_biwt = (~ core_wten) & cfg_mul_bypass_rsc_triosy_obj_iswt0;
  assign cfg_mul_bypass_rsc_triosy_obj_bdwt = cfg_mul_bypass_rsc_triosy_obj_oswt
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_out_rsci_oswt, chn_mul_out_rsci_bawt,
      chn_mul_out_rsci_wen_comp, chn_mul_out_rsci_biwt, chn_mul_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_out_rsci_oswt;
  output chn_mul_out_rsci_bawt;
  output chn_mul_out_rsci_wen_comp;
  input chn_mul_out_rsci_biwt;
  input chn_mul_out_rsci_bdwt;


  // Interconnect Declarations
  reg chn_mul_out_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_mul_out_rsci_bawt = chn_mul_out_rsci_biwt | chn_mul_out_rsci_bcwt;
  assign chn_mul_out_rsci_wen_comp = (~ chn_mul_out_rsci_oswt) | chn_mul_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_mul_out_rsci_bcwt <= ~((~(chn_mul_out_rsci_bcwt | chn_mul_out_rsci_biwt))
          | chn_mul_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_out_rsci_oswt, core_wen, core_wten, chn_mul_out_rsci_iswt0,
      chn_mul_out_rsci_ld_core_psct, chn_mul_out_rsci_biwt, chn_mul_out_rsci_bdwt,
      chn_mul_out_rsci_ld_core_sct, chn_mul_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_out_rsci_iswt0;
  input chn_mul_out_rsci_ld_core_psct;
  output chn_mul_out_rsci_biwt;
  output chn_mul_out_rsci_bdwt;
  output chn_mul_out_rsci_ld_core_sct;
  input chn_mul_out_rsci_vd;


  // Interconnect Declarations
  wire chn_mul_out_rsci_ogwt;
  wire chn_mul_out_rsci_pdswt0;
  reg chn_mul_out_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_mul_out_rsci_pdswt0 = (~ core_wten) & chn_mul_out_rsci_iswt0;
  assign chn_mul_out_rsci_biwt = chn_mul_out_rsci_ogwt & chn_mul_out_rsci_vd;
  assign chn_mul_out_rsci_ogwt = chn_mul_out_rsci_pdswt0 | chn_mul_out_rsci_icwt;
  assign chn_mul_out_rsci_bdwt = chn_mul_out_rsci_oswt & core_wen;
  assign chn_mul_out_rsci_ld_core_sct = chn_mul_out_rsci_ld_core_psct & chn_mul_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_mul_out_rsci_icwt <= ~((~(chn_mul_out_rsci_icwt | chn_mul_out_rsci_pdswt0))
          | chn_mul_out_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_op_rsci_oswt, chn_mul_op_rsci_bawt, chn_mul_op_rsci_wen_comp,
      chn_mul_op_rsci_d_mxwt, chn_mul_op_rsci_biwt, chn_mul_op_rsci_bdwt, chn_mul_op_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_op_rsci_oswt;
  output chn_mul_op_rsci_bawt;
  output chn_mul_op_rsci_wen_comp;
  output [127:0] chn_mul_op_rsci_d_mxwt;
  input chn_mul_op_rsci_biwt;
  input chn_mul_op_rsci_bdwt;
  input [127:0] chn_mul_op_rsci_d;


  // Interconnect Declarations
  reg chn_mul_op_rsci_bcwt;
  reg [127:0] chn_mul_op_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_mul_op_rsci_bawt = chn_mul_op_rsci_biwt | chn_mul_op_rsci_bcwt;
  assign chn_mul_op_rsci_wen_comp = (~ chn_mul_op_rsci_oswt) | chn_mul_op_rsci_bawt;
  assign chn_mul_op_rsci_d_mxwt = MUX_v_128_2_2(chn_mul_op_rsci_d, chn_mul_op_rsci_d_bfwt,
      chn_mul_op_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_op_rsci_bcwt <= 1'b0;
      chn_mul_op_rsci_d_bfwt <= 128'b0;
    end
    else begin
      chn_mul_op_rsci_bcwt <= ~((~(chn_mul_op_rsci_bcwt | chn_mul_op_rsci_biwt))
          | chn_mul_op_rsci_bdwt);
      chn_mul_op_rsci_d_bfwt <= chn_mul_op_rsci_d_mxwt;
    end
  end

  function [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_op_rsci_oswt, core_wen, core_wten, chn_mul_op_rsci_iswt0,
      chn_mul_op_rsci_ld_core_psct, chn_mul_op_rsci_biwt, chn_mul_op_rsci_bdwt, chn_mul_op_rsci_ld_core_sct,
      chn_mul_op_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_op_rsci_iswt0;
  input chn_mul_op_rsci_ld_core_psct;
  output chn_mul_op_rsci_biwt;
  output chn_mul_op_rsci_bdwt;
  output chn_mul_op_rsci_ld_core_sct;
  input chn_mul_op_rsci_vd;


  // Interconnect Declarations
  wire chn_mul_op_rsci_ogwt;
  wire chn_mul_op_rsci_pdswt0;
  reg chn_mul_op_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_mul_op_rsci_pdswt0 = (~ core_wten) & chn_mul_op_rsci_iswt0;
  assign chn_mul_op_rsci_biwt = chn_mul_op_rsci_ogwt & chn_mul_op_rsci_vd;
  assign chn_mul_op_rsci_ogwt = chn_mul_op_rsci_pdswt0 | chn_mul_op_rsci_icwt;
  assign chn_mul_op_rsci_bdwt = chn_mul_op_rsci_oswt & core_wen;
  assign chn_mul_op_rsci_ld_core_sct = chn_mul_op_rsci_ld_core_psct & chn_mul_op_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_op_rsci_icwt <= 1'b0;
    end
    else begin
      chn_mul_op_rsci_icwt <= ~((~(chn_mul_op_rsci_icwt | chn_mul_op_rsci_pdswt0))
          | chn_mul_op_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsci_oswt, chn_mul_in_rsci_bawt, chn_mul_in_rsci_wen_comp,
      chn_mul_in_rsci_d_mxwt, chn_mul_in_rsci_biwt, chn_mul_in_rsci_bdwt, chn_mul_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_in_rsci_oswt;
  output chn_mul_in_rsci_bawt;
  output chn_mul_in_rsci_wen_comp;
  output [127:0] chn_mul_in_rsci_d_mxwt;
  input chn_mul_in_rsci_biwt;
  input chn_mul_in_rsci_bdwt;
  input [127:0] chn_mul_in_rsci_d;


  // Interconnect Declarations
  reg chn_mul_in_rsci_bcwt;
  reg [127:0] chn_mul_in_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_mul_in_rsci_bawt = chn_mul_in_rsci_biwt | chn_mul_in_rsci_bcwt;
  assign chn_mul_in_rsci_wen_comp = (~ chn_mul_in_rsci_oswt) | chn_mul_in_rsci_bawt;
  assign chn_mul_in_rsci_d_mxwt = MUX_v_128_2_2(chn_mul_in_rsci_d, chn_mul_in_rsci_d_bfwt,
      chn_mul_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_bcwt <= 1'b0;
      chn_mul_in_rsci_d_bfwt <= 128'b0;
    end
    else begin
      chn_mul_in_rsci_bcwt <= ~((~(chn_mul_in_rsci_bcwt | chn_mul_in_rsci_biwt))
          | chn_mul_in_rsci_bdwt);
      chn_mul_in_rsci_d_bfwt <= chn_mul_in_rsci_d_mxwt;
    end
  end

  function [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsci_oswt, core_wen, chn_mul_in_rsci_iswt0,
      chn_mul_in_rsci_ld_core_psct, core_wten, chn_mul_in_rsci_biwt, chn_mul_in_rsci_bdwt,
      chn_mul_in_rsci_ld_core_sct, chn_mul_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_mul_in_rsci_oswt;
  input core_wen;
  input chn_mul_in_rsci_iswt0;
  input chn_mul_in_rsci_ld_core_psct;
  input core_wten;
  output chn_mul_in_rsci_biwt;
  output chn_mul_in_rsci_bdwt;
  output chn_mul_in_rsci_ld_core_sct;
  input chn_mul_in_rsci_vd;


  // Interconnect Declarations
  wire chn_mul_in_rsci_ogwt;
  wire chn_mul_in_rsci_pdswt0;
  reg chn_mul_in_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_mul_in_rsci_pdswt0 = (~ core_wten) & chn_mul_in_rsci_iswt0;
  assign chn_mul_in_rsci_biwt = chn_mul_in_rsci_ogwt & chn_mul_in_rsci_vd;
  assign chn_mul_in_rsci_ogwt = chn_mul_in_rsci_pdswt0 | chn_mul_in_rsci_icwt;
  assign chn_mul_in_rsci_bdwt = chn_mul_in_rsci_oswt & core_wen;
  assign chn_mul_in_rsci_ld_core_sct = chn_mul_in_rsci_ld_core_psct & chn_mul_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_mul_in_rsci_icwt <= ~((~(chn_mul_in_rsci_icwt | chn_mul_in_rsci_pdswt0))
          | chn_mul_in_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_alu_algo_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_alu_algo_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_alu_op_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_alu_op_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_alu_src_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_alu_src_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_cfg_alu_bypass_rsc_triosy_obj_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_cfg_alu_bypass_rsc_triosy_obj_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_chn_alu_out_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_chn_alu_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_chn_alu_op_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_chn_alu_op_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_chn_alu_in_rsci_unreg
// ------------------------------------------------------------------


module SDP_Y_CORE_chn_alu_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for Y_alu_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : Y_alu_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_staller
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_alu_in_rsci_wen_comp, core_wten,
      chn_alu_op_rsci_wen_comp, chn_alu_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_alu_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_alu_op_rsci_wen_comp;
  input chn_alu_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_alu_in_rsci_wen_comp & chn_alu_op_rsci_wen_comp & chn_alu_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_algo_rsc_triosy_obj_bawt, cfg_alu_algo_rsc_triosy_obj_biwt,
      cfg_alu_algo_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_algo_rsc_triosy_obj_bawt;
  input cfg_alu_algo_rsc_triosy_obj_biwt;
  input cfg_alu_algo_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_alu_algo_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_algo_rsc_triosy_obj_bawt = cfg_alu_algo_rsc_triosy_obj_biwt | cfg_alu_algo_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_algo_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_algo_rsc_triosy_obj_bcwt |
          cfg_alu_algo_rsc_triosy_obj_biwt)) | cfg_alu_algo_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl (
  cfg_alu_algo_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_algo_rsc_triosy_obj_iswt0,
      cfg_alu_algo_rsc_triosy_obj_biwt, cfg_alu_algo_rsc_triosy_obj_bdwt
);
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_algo_rsc_triosy_obj_iswt0;
  output cfg_alu_algo_rsc_triosy_obj_biwt;
  output cfg_alu_algo_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_algo_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_algo_rsc_triosy_obj_iswt0;
  assign cfg_alu_algo_rsc_triosy_obj_bdwt = cfg_alu_algo_rsc_triosy_obj_oswt & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_op_rsc_triosy_obj_bawt, cfg_alu_op_rsc_triosy_obj_biwt,
      cfg_alu_op_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_op_rsc_triosy_obj_bawt;
  input cfg_alu_op_rsc_triosy_obj_biwt;
  input cfg_alu_op_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_alu_op_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_op_rsc_triosy_obj_bawt = cfg_alu_op_rsc_triosy_obj_biwt | cfg_alu_op_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_op_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_op_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_op_rsc_triosy_obj_bcwt | cfg_alu_op_rsc_triosy_obj_biwt))
          | cfg_alu_op_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl (
  cfg_alu_op_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_op_rsc_triosy_obj_iswt0,
      cfg_alu_op_rsc_triosy_obj_biwt, cfg_alu_op_rsc_triosy_obj_bdwt
);
  input cfg_alu_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_op_rsc_triosy_obj_iswt0;
  output cfg_alu_op_rsc_triosy_obj_biwt;
  output cfg_alu_op_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_op_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_op_rsc_triosy_obj_iswt0;
  assign cfg_alu_op_rsc_triosy_obj_bdwt = cfg_alu_op_rsc_triosy_obj_oswt & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_src_rsc_triosy_obj_bawt, cfg_alu_src_rsc_triosy_obj_biwt,
      cfg_alu_src_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_src_rsc_triosy_obj_bawt;
  input cfg_alu_src_rsc_triosy_obj_biwt;
  input cfg_alu_src_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_alu_src_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_src_rsc_triosy_obj_bawt = cfg_alu_src_rsc_triosy_obj_biwt | cfg_alu_src_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_src_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_src_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_src_rsc_triosy_obj_bcwt | cfg_alu_src_rsc_triosy_obj_biwt))
          | cfg_alu_src_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl (
  cfg_alu_src_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_src_rsc_triosy_obj_iswt0,
      cfg_alu_src_rsc_triosy_obj_biwt, cfg_alu_src_rsc_triosy_obj_bdwt
);
  input cfg_alu_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_src_rsc_triosy_obj_iswt0;
  output cfg_alu_src_rsc_triosy_obj_biwt;
  output cfg_alu_src_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_src_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_src_rsc_triosy_obj_iswt0;
  assign cfg_alu_src_rsc_triosy_obj_bdwt = cfg_alu_src_rsc_triosy_obj_oswt & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp
    (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_bypass_rsc_triosy_obj_bawt, cfg_alu_bypass_rsc_triosy_obj_biwt,
      cfg_alu_bypass_rsc_triosy_obj_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_bypass_rsc_triosy_obj_bawt;
  input cfg_alu_bypass_rsc_triosy_obj_biwt;
  input cfg_alu_bypass_rsc_triosy_obj_bdwt;


  // Interconnect Declarations
  reg cfg_alu_bypass_rsc_triosy_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_bypass_rsc_triosy_obj_bawt = cfg_alu_bypass_rsc_triosy_obj_biwt
      | cfg_alu_bypass_rsc_triosy_obj_bcwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_bypass_rsc_triosy_obj_bcwt <= 1'b0;
    end
    else begin
      cfg_alu_bypass_rsc_triosy_obj_bcwt <= ~((~(cfg_alu_bypass_rsc_triosy_obj_bcwt
          | cfg_alu_bypass_rsc_triosy_obj_biwt)) | cfg_alu_bypass_rsc_triosy_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl
    (
  cfg_alu_bypass_rsc_triosy_obj_oswt, core_wen, core_wten, cfg_alu_bypass_rsc_triosy_obj_iswt0,
      cfg_alu_bypass_rsc_triosy_obj_biwt, cfg_alu_bypass_rsc_triosy_obj_bdwt
);
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_bypass_rsc_triosy_obj_iswt0;
  output cfg_alu_bypass_rsc_triosy_obj_biwt;
  output cfg_alu_bypass_rsc_triosy_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign cfg_alu_bypass_rsc_triosy_obj_biwt = (~ core_wten) & cfg_alu_bypass_rsc_triosy_obj_iswt0;
  assign cfg_alu_bypass_rsc_triosy_obj_bdwt = cfg_alu_bypass_rsc_triosy_obj_oswt
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_out_rsci_oswt, chn_alu_out_rsci_bawt,
      chn_alu_out_rsci_wen_comp, chn_alu_out_rsci_biwt, chn_alu_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_out_rsci_oswt;
  output chn_alu_out_rsci_bawt;
  output chn_alu_out_rsci_wen_comp;
  input chn_alu_out_rsci_biwt;
  input chn_alu_out_rsci_bdwt;


  // Interconnect Declarations
  reg chn_alu_out_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_alu_out_rsci_bawt = chn_alu_out_rsci_biwt | chn_alu_out_rsci_bcwt;
  assign chn_alu_out_rsci_wen_comp = (~ chn_alu_out_rsci_oswt) | chn_alu_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_alu_out_rsci_bcwt <= ~((~(chn_alu_out_rsci_bcwt | chn_alu_out_rsci_biwt))
          | chn_alu_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_out_rsci_oswt, core_wen, core_wten, chn_alu_out_rsci_iswt0,
      chn_alu_out_rsci_ld_core_psct, chn_alu_out_rsci_biwt, chn_alu_out_rsci_bdwt,
      chn_alu_out_rsci_ld_core_sct, chn_alu_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_out_rsci_iswt0;
  input chn_alu_out_rsci_ld_core_psct;
  output chn_alu_out_rsci_biwt;
  output chn_alu_out_rsci_bdwt;
  output chn_alu_out_rsci_ld_core_sct;
  input chn_alu_out_rsci_vd;


  // Interconnect Declarations
  wire chn_alu_out_rsci_ogwt;
  wire chn_alu_out_rsci_pdswt0;
  reg chn_alu_out_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_alu_out_rsci_pdswt0 = (~ core_wten) & chn_alu_out_rsci_iswt0;
  assign chn_alu_out_rsci_biwt = chn_alu_out_rsci_ogwt & chn_alu_out_rsci_vd;
  assign chn_alu_out_rsci_ogwt = chn_alu_out_rsci_pdswt0 | chn_alu_out_rsci_icwt;
  assign chn_alu_out_rsci_bdwt = chn_alu_out_rsci_oswt & core_wen;
  assign chn_alu_out_rsci_ld_core_sct = chn_alu_out_rsci_ld_core_psct & chn_alu_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_alu_out_rsci_icwt <= ~((~(chn_alu_out_rsci_icwt | chn_alu_out_rsci_pdswt0))
          | chn_alu_out_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_op_rsci_oswt, chn_alu_op_rsci_bawt, chn_alu_op_rsci_wen_comp,
      chn_alu_op_rsci_d_mxwt, chn_alu_op_rsci_biwt, chn_alu_op_rsci_bdwt, chn_alu_op_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_op_rsci_oswt;
  output chn_alu_op_rsci_bawt;
  output chn_alu_op_rsci_wen_comp;
  output [127:0] chn_alu_op_rsci_d_mxwt;
  input chn_alu_op_rsci_biwt;
  input chn_alu_op_rsci_bdwt;
  input [127:0] chn_alu_op_rsci_d;


  // Interconnect Declarations
  reg chn_alu_op_rsci_bcwt;
  reg [127:0] chn_alu_op_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_alu_op_rsci_bawt = chn_alu_op_rsci_biwt | chn_alu_op_rsci_bcwt;
  assign chn_alu_op_rsci_wen_comp = (~ chn_alu_op_rsci_oswt) | chn_alu_op_rsci_bawt;
  assign chn_alu_op_rsci_d_mxwt = MUX_v_128_2_2(chn_alu_op_rsci_d, chn_alu_op_rsci_d_bfwt,
      chn_alu_op_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_op_rsci_bcwt <= 1'b0;
      chn_alu_op_rsci_d_bfwt <= 128'b0;
    end
    else begin
      chn_alu_op_rsci_bcwt <= ~((~(chn_alu_op_rsci_bcwt | chn_alu_op_rsci_biwt))
          | chn_alu_op_rsci_bdwt);
      chn_alu_op_rsci_d_bfwt <= chn_alu_op_rsci_d_mxwt;
    end
  end

  function [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_op_rsci_oswt, core_wen, core_wten, chn_alu_op_rsci_iswt0,
      chn_alu_op_rsci_ld_core_psct, chn_alu_op_rsci_biwt, chn_alu_op_rsci_bdwt, chn_alu_op_rsci_ld_core_sct,
      chn_alu_op_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_op_rsci_iswt0;
  input chn_alu_op_rsci_ld_core_psct;
  output chn_alu_op_rsci_biwt;
  output chn_alu_op_rsci_bdwt;
  output chn_alu_op_rsci_ld_core_sct;
  input chn_alu_op_rsci_vd;


  // Interconnect Declarations
  wire chn_alu_op_rsci_ogwt;
  wire chn_alu_op_rsci_pdswt0;
  reg chn_alu_op_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_alu_op_rsci_pdswt0 = (~ core_wten) & chn_alu_op_rsci_iswt0;
  assign chn_alu_op_rsci_biwt = chn_alu_op_rsci_ogwt & chn_alu_op_rsci_vd;
  assign chn_alu_op_rsci_ogwt = chn_alu_op_rsci_pdswt0 | chn_alu_op_rsci_icwt;
  assign chn_alu_op_rsci_bdwt = chn_alu_op_rsci_oswt & core_wen;
  assign chn_alu_op_rsci_ld_core_sct = chn_alu_op_rsci_ld_core_psct & chn_alu_op_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_op_rsci_icwt <= 1'b0;
    end
    else begin
      chn_alu_op_rsci_icwt <= ~((~(chn_alu_op_rsci_icwt | chn_alu_op_rsci_pdswt0))
          | chn_alu_op_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsci_oswt, chn_alu_in_rsci_bawt, chn_alu_in_rsci_wen_comp,
      chn_alu_in_rsci_d_mxwt, chn_alu_in_rsci_biwt, chn_alu_in_rsci_bdwt, chn_alu_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_in_rsci_oswt;
  output chn_alu_in_rsci_bawt;
  output chn_alu_in_rsci_wen_comp;
  output [127:0] chn_alu_in_rsci_d_mxwt;
  input chn_alu_in_rsci_biwt;
  input chn_alu_in_rsci_bdwt;
  input [127:0] chn_alu_in_rsci_d;


  // Interconnect Declarations
  reg chn_alu_in_rsci_bcwt;
  reg [127:0] chn_alu_in_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_alu_in_rsci_bawt = chn_alu_in_rsci_biwt | chn_alu_in_rsci_bcwt;
  assign chn_alu_in_rsci_wen_comp = (~ chn_alu_in_rsci_oswt) | chn_alu_in_rsci_bawt;
  assign chn_alu_in_rsci_d_mxwt = MUX_v_128_2_2(chn_alu_in_rsci_d, chn_alu_in_rsci_d_bfwt,
      chn_alu_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_bcwt <= 1'b0;
      chn_alu_in_rsci_d_bfwt <= 128'b0;
    end
    else begin
      chn_alu_in_rsci_bcwt <= ~((~(chn_alu_in_rsci_bcwt | chn_alu_in_rsci_biwt))
          | chn_alu_in_rsci_bdwt);
      chn_alu_in_rsci_d_bfwt <= chn_alu_in_rsci_d_mxwt;
    end
  end

  function [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsci_oswt, core_wen, chn_alu_in_rsci_iswt0,
      chn_alu_in_rsci_ld_core_psct, core_wten, chn_alu_in_rsci_biwt, chn_alu_in_rsci_bdwt,
      chn_alu_in_rsci_ld_core_sct, chn_alu_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_alu_in_rsci_oswt;
  input core_wen;
  input chn_alu_in_rsci_iswt0;
  input chn_alu_in_rsci_ld_core_psct;
  input core_wten;
  output chn_alu_in_rsci_biwt;
  output chn_alu_in_rsci_bdwt;
  output chn_alu_in_rsci_ld_core_sct;
  input chn_alu_in_rsci_vd;


  // Interconnect Declarations
  wire chn_alu_in_rsci_ogwt;
  wire chn_alu_in_rsci_pdswt0;
  reg chn_alu_in_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_alu_in_rsci_pdswt0 = (~ core_wten) & chn_alu_in_rsci_iswt0;
  assign chn_alu_in_rsci_biwt = chn_alu_in_rsci_ogwt & chn_alu_in_rsci_vd;
  assign chn_alu_in_rsci_ogwt = chn_alu_in_rsci_pdswt0 | chn_alu_in_rsci_icwt;
  assign chn_alu_in_rsci_bdwt = chn_alu_in_rsci_oswt & core_wen;
  assign chn_alu_in_rsci_ld_core_sct = chn_alu_in_rsci_ld_core_psct & chn_alu_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_alu_in_rsci_icwt <= ~((~(chn_alu_in_rsci_icwt | chn_alu_in_rsci_pdswt0))
          | chn_alu_in_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_truncate_rsc_triosy_lz, cfg_truncate_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_truncate_rsc_triosy_obj_iswt0, cfg_truncate_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_truncate_rsc_triosy_lz;
  input cfg_truncate_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_truncate_rsc_triosy_obj_iswt0;
  output cfg_truncate_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_truncate_rsc_triosy_obj_biwt;
  wire cfg_truncate_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_truncate_rsc_triosy_obj (
      .ld(cfg_truncate_rsc_triosy_obj_biwt),
      .lz(cfg_truncate_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_ctrl Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_ctrl_inst
      (
      .cfg_truncate_rsc_triosy_obj_oswt(cfg_truncate_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_truncate_rsc_triosy_obj_iswt0(cfg_truncate_rsc_triosy_obj_iswt0),
      .cfg_truncate_rsc_triosy_obj_biwt(cfg_truncate_rsc_triosy_obj_biwt),
      .cfg_truncate_rsc_triosy_obj_bdwt(cfg_truncate_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_dp Y_mul_core_cfg_truncate_rsc_triosy_obj_cfg_truncate_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_truncate_rsc_triosy_obj_bawt(cfg_truncate_rsc_triosy_obj_bawt),
      .cfg_truncate_rsc_triosy_obj_biwt(cfg_truncate_rsc_triosy_obj_biwt),
      .cfg_truncate_rsc_triosy_obj_bdwt(cfg_truncate_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_op_rsc_triosy_lz, cfg_mul_op_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_op_rsc_triosy_obj_iswt0, cfg_mul_op_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_op_rsc_triosy_lz;
  input cfg_mul_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_op_rsc_triosy_obj_iswt0;
  output cfg_mul_op_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_mul_op_rsc_triosy_obj_biwt;
  wire cfg_mul_op_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_op_rsc_triosy_obj (
      .ld(cfg_mul_op_rsc_triosy_obj_biwt),
      .lz(cfg_mul_op_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_op_rsc_triosy_obj_iswt0(cfg_mul_op_rsc_triosy_obj_iswt0),
      .cfg_mul_op_rsc_triosy_obj_biwt(cfg_mul_op_rsc_triosy_obj_biwt),
      .cfg_mul_op_rsc_triosy_obj_bdwt(cfg_mul_op_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp Y_mul_core_cfg_mul_op_rsc_triosy_obj_cfg_mul_op_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_op_rsc_triosy_obj_bawt(cfg_mul_op_rsc_triosy_obj_bawt),
      .cfg_mul_op_rsc_triosy_obj_biwt(cfg_mul_op_rsc_triosy_obj_biwt),
      .cfg_mul_op_rsc_triosy_obj_bdwt(cfg_mul_op_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_src_rsc_triosy_lz, cfg_mul_src_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_src_rsc_triosy_obj_iswt0, cfg_mul_src_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_src_rsc_triosy_lz;
  input cfg_mul_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_src_rsc_triosy_obj_iswt0;
  output cfg_mul_src_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_mul_src_rsc_triosy_obj_biwt;
  wire cfg_mul_src_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_src_rsc_triosy_obj (
      .ld(cfg_mul_src_rsc_triosy_obj_biwt),
      .lz(cfg_mul_src_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_src_rsc_triosy_obj_iswt0(cfg_mul_src_rsc_triosy_obj_iswt0),
      .cfg_mul_src_rsc_triosy_obj_biwt(cfg_mul_src_rsc_triosy_obj_biwt),
      .cfg_mul_src_rsc_triosy_obj_bdwt(cfg_mul_src_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp Y_mul_core_cfg_mul_src_rsc_triosy_obj_cfg_mul_src_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_src_rsc_triosy_obj_bawt(cfg_mul_src_rsc_triosy_obj_bawt),
      .cfg_mul_src_rsc_triosy_obj_biwt(cfg_mul_src_rsc_triosy_obj_biwt),
      .cfg_mul_src_rsc_triosy_obj_bdwt(cfg_mul_src_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_prelu_rsc_triosy_lz, cfg_mul_prelu_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_prelu_rsc_triosy_obj_iswt0, cfg_mul_prelu_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_prelu_rsc_triosy_lz;
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_prelu_rsc_triosy_obj_iswt0;
  output cfg_mul_prelu_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_mul_prelu_rsc_triosy_obj_biwt;
  wire cfg_mul_prelu_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_prelu_rsc_triosy_obj (
      .ld(cfg_mul_prelu_rsc_triosy_obj_biwt),
      .lz(cfg_mul_prelu_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_prelu_rsc_triosy_obj_iswt0(cfg_mul_prelu_rsc_triosy_obj_iswt0),
      .cfg_mul_prelu_rsc_triosy_obj_biwt(cfg_mul_prelu_rsc_triosy_obj_biwt),
      .cfg_mul_prelu_rsc_triosy_obj_bdwt(cfg_mul_prelu_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_cfg_mul_prelu_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_prelu_rsc_triosy_obj_bawt(cfg_mul_prelu_rsc_triosy_obj_bawt),
      .cfg_mul_prelu_rsc_triosy_obj_biwt(cfg_mul_prelu_rsc_triosy_obj_biwt),
      .cfg_mul_prelu_rsc_triosy_obj_bdwt(cfg_mul_prelu_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_mul_bypass_rsc_triosy_lz, cfg_mul_bypass_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_mul_bypass_rsc_triosy_obj_iswt0, cfg_mul_bypass_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_mul_bypass_rsc_triosy_lz;
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_mul_bypass_rsc_triosy_obj_iswt0;
  output cfg_mul_bypass_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_mul_bypass_rsc_triosy_obj_biwt;
  wire cfg_mul_bypass_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_mul_bypass_rsc_triosy_obj (
      .ld(cfg_mul_bypass_rsc_triosy_obj_biwt),
      .lz(cfg_mul_bypass_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_ctrl_inst
      (
      .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_bypass_rsc_triosy_obj_iswt0(cfg_mul_bypass_rsc_triosy_obj_iswt0),
      .cfg_mul_bypass_rsc_triosy_obj_biwt(cfg_mul_bypass_rsc_triosy_obj_biwt),
      .cfg_mul_bypass_rsc_triosy_obj_bdwt(cfg_mul_bypass_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_cfg_mul_bypass_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_bypass_rsc_triosy_obj_bawt(cfg_mul_bypass_rsc_triosy_obj_bawt),
      .cfg_mul_bypass_rsc_triosy_obj_biwt(cfg_mul_bypass_rsc_triosy_obj_biwt),
      .cfg_mul_bypass_rsc_triosy_obj_bdwt(cfg_mul_bypass_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_out_rsc_z, chn_mul_out_rsc_vz, chn_mul_out_rsc_lz,
      chn_mul_out_rsci_oswt, core_wen, core_wten, chn_mul_out_rsci_iswt0, chn_mul_out_rsci_bawt,
      chn_mul_out_rsci_wen_comp, chn_mul_out_rsci_ld_core_psct, chn_mul_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [127:0] chn_mul_out_rsc_z;
  input chn_mul_out_rsc_vz;
  output chn_mul_out_rsc_lz;
  input chn_mul_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_out_rsci_iswt0;
  output chn_mul_out_rsci_bawt;
  output chn_mul_out_rsci_wen_comp;
  input chn_mul_out_rsci_ld_core_psct;
  input [127:0] chn_mul_out_rsci_d;


  // Interconnect Declarations
  wire chn_mul_out_rsci_biwt;
  wire chn_mul_out_rsci_bdwt;
  wire chn_mul_out_rsci_ld_core_sct;
  wire chn_mul_out_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_out_stdreg_wait_v1 #(.rscid(32'sd9),
  .width(32'sd128)) chn_mul_out_rsci (
      .ld(chn_mul_out_rsci_ld_core_sct),
      .vd(chn_mul_out_rsci_vd),
      .d(chn_mul_out_rsci_d),
      .lz(chn_mul_out_rsc_lz),
      .vz(chn_mul_out_rsc_vz),
      .z(chn_mul_out_rsc_z)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_out_rsci_iswt0(chn_mul_out_rsci_iswt0),
      .chn_mul_out_rsci_ld_core_psct(chn_mul_out_rsci_ld_core_psct),
      .chn_mul_out_rsci_biwt(chn_mul_out_rsci_biwt),
      .chn_mul_out_rsci_bdwt(chn_mul_out_rsci_bdwt),
      .chn_mul_out_rsci_ld_core_sct(chn_mul_out_rsci_ld_core_sct),
      .chn_mul_out_rsci_vd(chn_mul_out_rsci_vd)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp Y_mul_core_chn_mul_out_rsci_chn_mul_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .chn_mul_out_rsci_bawt(chn_mul_out_rsci_bawt),
      .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp),
      .chn_mul_out_rsci_biwt(chn_mul_out_rsci_biwt),
      .chn_mul_out_rsci_bdwt(chn_mul_out_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_op_rsc_z, chn_mul_op_rsc_vz, chn_mul_op_rsc_lz,
      chn_mul_op_rsci_oswt, core_wen, core_wten, chn_mul_op_rsci_iswt0, chn_mul_op_rsci_bawt,
      chn_mul_op_rsci_wen_comp, chn_mul_op_rsci_ld_core_psct, chn_mul_op_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  input chn_mul_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_mul_op_rsci_iswt0;
  output chn_mul_op_rsci_bawt;
  output chn_mul_op_rsci_wen_comp;
  input chn_mul_op_rsci_ld_core_psct;
  output [127:0] chn_mul_op_rsci_d_mxwt;


  // Interconnect Declarations
  wire chn_mul_op_rsci_biwt;
  wire chn_mul_op_rsci_bdwt;
  wire chn_mul_op_rsci_ld_core_sct;
  wire chn_mul_op_rsci_vd;
  wire [127:0] chn_mul_op_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_in_wire_wait_v1 #(.rscid(32'sd2),
  .width(32'sd128)) chn_mul_op_rsci (
      .ld(chn_mul_op_rsci_ld_core_sct),
      .vd(chn_mul_op_rsci_vd),
      .d(chn_mul_op_rsci_d),
      .lz(chn_mul_op_rsc_lz),
      .vz(chn_mul_op_rsc_vz),
      .z(chn_mul_op_rsc_z)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_op_rsci_iswt0(chn_mul_op_rsci_iswt0),
      .chn_mul_op_rsci_ld_core_psct(chn_mul_op_rsci_ld_core_psct),
      .chn_mul_op_rsci_biwt(chn_mul_op_rsci_biwt),
      .chn_mul_op_rsci_bdwt(chn_mul_op_rsci_bdwt),
      .chn_mul_op_rsci_ld_core_sct(chn_mul_op_rsci_ld_core_sct),
      .chn_mul_op_rsci_vd(chn_mul_op_rsci_vd)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp Y_mul_core_chn_mul_op_rsci_chn_mul_op_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .chn_mul_op_rsci_bawt(chn_mul_op_rsci_bawt),
      .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
      .chn_mul_op_rsci_d_mxwt(chn_mul_op_rsci_d_mxwt),
      .chn_mul_op_rsci_biwt(chn_mul_op_rsci_biwt),
      .chn_mul_op_rsci_bdwt(chn_mul_op_rsci_bdwt),
      .chn_mul_op_rsci_d(chn_mul_op_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_z, chn_mul_in_rsc_vz, chn_mul_in_rsc_lz,
      chn_mul_in_rsci_oswt, core_wen, chn_mul_in_rsci_iswt0, chn_mul_in_rsci_bawt,
      chn_mul_in_rsci_wen_comp, chn_mul_in_rsci_ld_core_psct, chn_mul_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_mul_in_rsc_z;
  input chn_mul_in_rsc_vz;
  output chn_mul_in_rsc_lz;
  input chn_mul_in_rsci_oswt;
  input core_wen;
  input chn_mul_in_rsci_iswt0;
  output chn_mul_in_rsci_bawt;
  output chn_mul_in_rsci_wen_comp;
  input chn_mul_in_rsci_ld_core_psct;
  output [127:0] chn_mul_in_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_mul_in_rsci_biwt;
  wire chn_mul_in_rsci_bdwt;
  wire chn_mul_in_rsci_ld_core_sct;
  wire chn_mul_in_rsci_vd;
  wire [127:0] chn_mul_in_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd128)) chn_mul_in_rsci (
      .ld(chn_mul_in_rsci_ld_core_sct),
      .vd(chn_mul_in_rsci_vd),
      .d(chn_mul_in_rsci_d),
      .lz(chn_mul_in_rsc_lz),
      .vz(chn_mul_in_rsc_vz),
      .z(chn_mul_in_rsc_z)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_mul_in_rsci_iswt0(chn_mul_in_rsci_iswt0),
      .chn_mul_in_rsci_ld_core_psct(chn_mul_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_mul_in_rsci_biwt(chn_mul_in_rsci_biwt),
      .chn_mul_in_rsci_bdwt(chn_mul_in_rsci_bdwt),
      .chn_mul_in_rsci_ld_core_sct(chn_mul_in_rsci_ld_core_sct),
      .chn_mul_in_rsci_vd(chn_mul_in_rsci_vd)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp Y_mul_core_chn_mul_in_rsci_chn_mul_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .chn_mul_in_rsci_bawt(chn_mul_in_rsci_bawt),
      .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
      .chn_mul_in_rsci_d_mxwt(chn_mul_in_rsci_d_mxwt),
      .chn_mul_in_rsci_biwt(chn_mul_in_rsci_biwt),
      .chn_mul_in_rsci_bdwt(chn_mul_in_rsci_bdwt),
      .chn_mul_in_rsci_d(chn_mul_in_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_algo_rsc_triosy_lz, cfg_alu_algo_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_algo_rsc_triosy_obj_iswt0, cfg_alu_algo_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_algo_rsc_triosy_lz;
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_algo_rsc_triosy_obj_iswt0;
  output cfg_alu_algo_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_alu_algo_rsc_triosy_obj_biwt;
  wire cfg_alu_algo_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_algo_rsc_triosy_obj (
      .ld(cfg_alu_algo_rsc_triosy_obj_biwt),
      .lz(cfg_alu_algo_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_algo_rsc_triosy_obj_iswt0(cfg_alu_algo_rsc_triosy_obj_iswt0),
      .cfg_alu_algo_rsc_triosy_obj_biwt(cfg_alu_algo_rsc_triosy_obj_biwt),
      .cfg_alu_algo_rsc_triosy_obj_bdwt(cfg_alu_algo_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp Y_alu_core_cfg_alu_algo_rsc_triosy_obj_cfg_alu_algo_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_algo_rsc_triosy_obj_bawt(cfg_alu_algo_rsc_triosy_obj_bawt),
      .cfg_alu_algo_rsc_triosy_obj_biwt(cfg_alu_algo_rsc_triosy_obj_biwt),
      .cfg_alu_algo_rsc_triosy_obj_bdwt(cfg_alu_algo_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_op_rsc_triosy_lz, cfg_alu_op_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_op_rsc_triosy_obj_iswt0, cfg_alu_op_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_op_rsc_triosy_lz;
  input cfg_alu_op_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_op_rsc_triosy_obj_iswt0;
  output cfg_alu_op_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_alu_op_rsc_triosy_obj_biwt;
  wire cfg_alu_op_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_op_rsc_triosy_obj (
      .ld(cfg_alu_op_rsc_triosy_obj_biwt),
      .lz(cfg_alu_op_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_op_rsc_triosy_obj_iswt0(cfg_alu_op_rsc_triosy_obj_iswt0),
      .cfg_alu_op_rsc_triosy_obj_biwt(cfg_alu_op_rsc_triosy_obj_biwt),
      .cfg_alu_op_rsc_triosy_obj_bdwt(cfg_alu_op_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp Y_alu_core_cfg_alu_op_rsc_triosy_obj_cfg_alu_op_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_op_rsc_triosy_obj_bawt(cfg_alu_op_rsc_triosy_obj_bawt),
      .cfg_alu_op_rsc_triosy_obj_biwt(cfg_alu_op_rsc_triosy_obj_biwt),
      .cfg_alu_op_rsc_triosy_obj_bdwt(cfg_alu_op_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_src_rsc_triosy_lz, cfg_alu_src_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_src_rsc_triosy_obj_iswt0, cfg_alu_src_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_src_rsc_triosy_lz;
  input cfg_alu_src_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_src_rsc_triosy_obj_iswt0;
  output cfg_alu_src_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_alu_src_rsc_triosy_obj_biwt;
  wire cfg_alu_src_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_src_rsc_triosy_obj (
      .ld(cfg_alu_src_rsc_triosy_obj_biwt),
      .lz(cfg_alu_src_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_src_rsc_triosy_obj_iswt0(cfg_alu_src_rsc_triosy_obj_iswt0),
      .cfg_alu_src_rsc_triosy_obj_biwt(cfg_alu_src_rsc_triosy_obj_biwt),
      .cfg_alu_src_rsc_triosy_obj_bdwt(cfg_alu_src_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp Y_alu_core_cfg_alu_src_rsc_triosy_obj_cfg_alu_src_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_src_rsc_triosy_obj_bawt(cfg_alu_src_rsc_triosy_obj_bawt),
      .cfg_alu_src_rsc_triosy_obj_biwt(cfg_alu_src_rsc_triosy_obj_biwt),
      .cfg_alu_src_rsc_triosy_obj_bdwt(cfg_alu_src_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj (
  nvdla_core_clk, nvdla_core_rstn, cfg_alu_bypass_rsc_triosy_lz, cfg_alu_bypass_rsc_triosy_obj_oswt,
      core_wen, core_wten, cfg_alu_bypass_rsc_triosy_obj_iswt0, cfg_alu_bypass_rsc_triosy_obj_bawt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output cfg_alu_bypass_rsc_triosy_lz;
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  input core_wen;
  input core_wten;
  input cfg_alu_bypass_rsc_triosy_obj_iswt0;
  output cfg_alu_bypass_rsc_triosy_obj_bawt;


  // Interconnect Declarations
  wire cfg_alu_bypass_rsc_triosy_obj_biwt;
  wire cfg_alu_bypass_rsc_triosy_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_io_sync_v1 #(.valid(32'sd0)) cfg_alu_bypass_rsc_triosy_obj (
      .ld(cfg_alu_bypass_rsc_triosy_obj_biwt),
      .lz(cfg_alu_bypass_rsc_triosy_lz)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_ctrl_inst
      (
      .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_bypass_rsc_triosy_obj_iswt0(cfg_alu_bypass_rsc_triosy_obj_iswt0),
      .cfg_alu_bypass_rsc_triosy_obj_biwt(cfg_alu_bypass_rsc_triosy_obj_biwt),
      .cfg_alu_bypass_rsc_triosy_obj_bdwt(cfg_alu_bypass_rsc_triosy_obj_bdwt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_cfg_alu_bypass_rsc_triosy_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_bypass_rsc_triosy_obj_bawt(cfg_alu_bypass_rsc_triosy_obj_bawt),
      .cfg_alu_bypass_rsc_triosy_obj_biwt(cfg_alu_bypass_rsc_triosy_obj_biwt),
      .cfg_alu_bypass_rsc_triosy_obj_bdwt(cfg_alu_bypass_rsc_triosy_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_out_rsc_z, chn_alu_out_rsc_vz, chn_alu_out_rsc_lz,
      chn_alu_out_rsci_oswt, core_wen, core_wten, chn_alu_out_rsci_iswt0, chn_alu_out_rsci_bawt,
      chn_alu_out_rsci_wen_comp, chn_alu_out_rsci_ld_core_psct, chn_alu_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [127:0] chn_alu_out_rsc_z;
  input chn_alu_out_rsc_vz;
  output chn_alu_out_rsc_lz;
  input chn_alu_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_out_rsci_iswt0;
  output chn_alu_out_rsci_bawt;
  output chn_alu_out_rsci_wen_comp;
  input chn_alu_out_rsci_ld_core_psct;
  input [127:0] chn_alu_out_rsci_d;


  // Interconnect Declarations
  wire chn_alu_out_rsci_biwt;
  wire chn_alu_out_rsci_bdwt;
  wire chn_alu_out_rsci_ld_core_sct;
  wire chn_alu_out_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_out_stdreg_wait_v1 #(.rscid(32'sd20),
  .width(32'sd128)) chn_alu_out_rsci (
      .ld(chn_alu_out_rsci_ld_core_sct),
      .vd(chn_alu_out_rsci_vd),
      .d(chn_alu_out_rsci_d),
      .lz(chn_alu_out_rsc_lz),
      .vz(chn_alu_out_rsc_vz),
      .z(chn_alu_out_rsc_z)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_out_rsci_iswt0(chn_alu_out_rsci_iswt0),
      .chn_alu_out_rsci_ld_core_psct(chn_alu_out_rsci_ld_core_psct),
      .chn_alu_out_rsci_biwt(chn_alu_out_rsci_biwt),
      .chn_alu_out_rsci_bdwt(chn_alu_out_rsci_bdwt),
      .chn_alu_out_rsci_ld_core_sct(chn_alu_out_rsci_ld_core_sct),
      .chn_alu_out_rsci_vd(chn_alu_out_rsci_vd)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp Y_alu_core_chn_alu_out_rsci_chn_alu_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .chn_alu_out_rsci_bawt(chn_alu_out_rsci_bawt),
      .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp),
      .chn_alu_out_rsci_biwt(chn_alu_out_rsci_biwt),
      .chn_alu_out_rsci_bdwt(chn_alu_out_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz,
      chn_alu_op_rsci_oswt, core_wen, core_wten, chn_alu_op_rsci_iswt0, chn_alu_op_rsci_bawt,
      chn_alu_op_rsci_wen_comp, chn_alu_op_rsci_ld_core_psct, chn_alu_op_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  input chn_alu_op_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_alu_op_rsci_iswt0;
  output chn_alu_op_rsci_bawt;
  output chn_alu_op_rsci_wen_comp;
  input chn_alu_op_rsci_ld_core_psct;
  output [127:0] chn_alu_op_rsci_d_mxwt;


  // Interconnect Declarations
  wire chn_alu_op_rsci_biwt;
  wire chn_alu_op_rsci_bdwt;
  wire chn_alu_op_rsci_ld_core_sct;
  wire chn_alu_op_rsci_vd;
  wire [127:0] chn_alu_op_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_in_wire_wait_v1 #(.rscid(32'sd14),
  .width(32'sd128)) chn_alu_op_rsci (
      .ld(chn_alu_op_rsci_ld_core_sct),
      .vd(chn_alu_op_rsci_vd),
      .d(chn_alu_op_rsci_d),
      .lz(chn_alu_op_rsc_lz),
      .vz(chn_alu_op_rsc_vz),
      .z(chn_alu_op_rsc_z)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_op_rsci_iswt0(chn_alu_op_rsci_iswt0),
      .chn_alu_op_rsci_ld_core_psct(chn_alu_op_rsci_ld_core_psct),
      .chn_alu_op_rsci_biwt(chn_alu_op_rsci_biwt),
      .chn_alu_op_rsci_bdwt(chn_alu_op_rsci_bdwt),
      .chn_alu_op_rsci_ld_core_sct(chn_alu_op_rsci_ld_core_sct),
      .chn_alu_op_rsci_vd(chn_alu_op_rsci_vd)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp Y_alu_core_chn_alu_op_rsci_chn_alu_op_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .chn_alu_op_rsci_bawt(chn_alu_op_rsci_bawt),
      .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
      .chn_alu_op_rsci_d_mxwt(chn_alu_op_rsci_d_mxwt),
      .chn_alu_op_rsci_biwt(chn_alu_op_rsci_biwt),
      .chn_alu_op_rsci_bdwt(chn_alu_op_rsci_bdwt),
      .chn_alu_op_rsci_d(chn_alu_op_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz,
      chn_alu_in_rsci_oswt, core_wen, chn_alu_in_rsci_iswt0, chn_alu_in_rsci_bawt,
      chn_alu_in_rsci_wen_comp, chn_alu_in_rsci_ld_core_psct, chn_alu_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_alu_in_rsc_z;
  input chn_alu_in_rsc_vz;
  output chn_alu_in_rsc_lz;
  input chn_alu_in_rsci_oswt;
  input core_wen;
  input chn_alu_in_rsci_iswt0;
  output chn_alu_in_rsci_bawt;
  output chn_alu_in_rsci_wen_comp;
  input chn_alu_in_rsci_ld_core_psct;
  output [127:0] chn_alu_in_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_alu_in_rsci_biwt;
  wire chn_alu_in_rsci_bdwt;
  wire chn_alu_in_rsci_ld_core_sct;
  wire chn_alu_in_rsci_vd;
  wire [127:0] chn_alu_in_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_in_wire_wait_v1 #(.rscid(32'sd13),
  .width(32'sd128)) chn_alu_in_rsci (
      .ld(chn_alu_in_rsci_ld_core_sct),
      .vd(chn_alu_in_rsci_vd),
      .d(chn_alu_in_rsci_d),
      .lz(chn_alu_in_rsc_lz),
      .vz(chn_alu_in_rsc_vz),
      .z(chn_alu_in_rsc_z)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_alu_in_rsci_iswt0(chn_alu_in_rsci_iswt0),
      .chn_alu_in_rsci_ld_core_psct(chn_alu_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_alu_in_rsci_biwt(chn_alu_in_rsci_biwt),
      .chn_alu_in_rsci_bdwt(chn_alu_in_rsci_bdwt),
      .chn_alu_in_rsci_ld_core_sct(chn_alu_in_rsci_ld_core_sct),
      .chn_alu_in_rsci_vd(chn_alu_in_rsci_vd)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp Y_alu_core_chn_alu_in_rsci_chn_alu_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .chn_alu_in_rsci_bawt(chn_alu_in_rsci_bawt),
      .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
      .chn_alu_in_rsci_d_mxwt(chn_alu_in_rsci_d_mxwt),
      .chn_alu_in_rsci_biwt(chn_alu_in_rsci_biwt),
      .chn_alu_in_rsci_bdwt(chn_alu_in_rsci_bdwt),
      .chn_alu_in_rsci_d(chn_alu_in_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul_core
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul_core (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_z, chn_mul_in_rsc_vz, chn_mul_in_rsc_lz,
      chn_mul_op_rsc_z, chn_mul_op_rsc_vz, chn_mul_op_rsc_lz, cfg_mul_bypass_rsc_triosy_lz,
      cfg_mul_prelu_rsc_triosy_lz, cfg_mul_src_rsc_triosy_lz, cfg_mul_op_rsc_triosy_lz,
      cfg_truncate_rsc_triosy_lz, cfg_precision, chn_mul_out_rsc_z, chn_mul_out_rsc_vz,
      chn_mul_out_rsc_lz, chn_mul_in_rsci_oswt, chn_mul_in_rsci_oswt_unreg, chn_mul_op_rsci_oswt,
      chn_mul_op_rsci_oswt_unreg, cfg_mul_bypass_rsci_d, cfg_mul_prelu_rsci_d, cfg_mul_src_rsci_d,
      cfg_mul_op_rsci_d, cfg_truncate_rsci_d, chn_mul_out_rsci_oswt, chn_mul_out_rsci_oswt_unreg,
      cfg_mul_bypass_rsc_triosy_obj_oswt, cfg_mul_prelu_rsc_triosy_obj_oswt, cfg_mul_src_rsc_triosy_obj_oswt,
      cfg_mul_op_rsc_triosy_obj_oswt, cfg_truncate_rsc_triosy_obj_oswt, cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_mul_in_rsc_z;
  input chn_mul_in_rsc_vz;
  output chn_mul_in_rsc_lz;
  input [127:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  output cfg_mul_bypass_rsc_triosy_lz;
  output cfg_mul_prelu_rsc_triosy_lz;
  output cfg_mul_src_rsc_triosy_lz;
  output cfg_mul_op_rsc_triosy_lz;
  output cfg_truncate_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [127:0] chn_mul_out_rsc_z;
  input chn_mul_out_rsc_vz;
  output chn_mul_out_rsc_lz;
  input chn_mul_in_rsci_oswt;
  output chn_mul_in_rsci_oswt_unreg;
  input chn_mul_op_rsci_oswt;
  output chn_mul_op_rsci_oswt_unreg;
  input cfg_mul_bypass_rsci_d;
  input cfg_mul_prelu_rsci_d;
  input cfg_mul_src_rsci_d;
  input [31:0] cfg_mul_op_rsci_d;
  input [9:0] cfg_truncate_rsci_d;
  input chn_mul_out_rsci_oswt;
  output chn_mul_out_rsci_oswt_unreg;
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  input cfg_mul_src_rsc_triosy_obj_oswt;
  input cfg_mul_op_rsc_triosy_obj_oswt;
  input cfg_truncate_rsc_triosy_obj_oswt;
  output cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff;


  // Interconnect Declarations
  wire core_wen;
  reg chn_mul_in_rsci_iswt0;
  wire chn_mul_in_rsci_bawt;
  wire chn_mul_in_rsci_wen_comp;
  reg chn_mul_in_rsci_ld_core_psct;
  wire [127:0] chn_mul_in_rsci_d_mxwt;
  wire core_wten;
  reg chn_mul_op_rsci_iswt0;
  wire chn_mul_op_rsci_bawt;
  wire chn_mul_op_rsci_wen_comp;
  reg chn_mul_op_rsci_ld_core_psct;
  wire [127:0] chn_mul_op_rsci_d_mxwt;
  reg chn_mul_out_rsci_iswt0;
  wire chn_mul_out_rsci_bawt;
  wire chn_mul_out_rsci_wen_comp;
  wire cfg_mul_bypass_rsc_triosy_obj_bawt;
  wire cfg_mul_prelu_rsc_triosy_obj_bawt;
  wire cfg_mul_src_rsc_triosy_obj_bawt;
  wire cfg_mul_op_rsc_triosy_obj_bawt;
  wire cfg_truncate_rsc_triosy_obj_bawt;
  reg chn_mul_out_rsci_d_127;
  reg [7:0] chn_mul_out_rsci_d_126_119;
  reg [21:0] chn_mul_out_rsci_d_118_97;
  reg chn_mul_out_rsci_d_96;
  reg chn_mul_out_rsci_d_95;
  reg [7:0] chn_mul_out_rsci_d_94_87;
  reg [21:0] chn_mul_out_rsci_d_86_65;
  reg chn_mul_out_rsci_d_64;
  reg chn_mul_out_rsci_d_63;
  reg [7:0] chn_mul_out_rsci_d_62_55;
  reg [21:0] chn_mul_out_rsci_d_54_33;
  reg chn_mul_out_rsci_d_32;
  reg chn_mul_out_rsci_d_31;
  reg [7:0] chn_mul_out_rsci_d_30_23;
  reg [21:0] chn_mul_out_rsci_d_22_1;
  reg chn_mul_out_rsci_d_0;
  wire [1:0] fsm_output;
  wire and_20_tmp;
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  wire and_18_tmp;
  wire [47:0] mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire [47:0] mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp;
  wire mul_mul_4_FpMantRNE_48U_24U_else_and_tmp;
  wire mul_mul_3_FpMantRNE_48U_24U_else_and_tmp;
  wire mul_mul_2_FpMantRNE_48U_24U_else_and_tmp;
  wire mul_mul_1_FpMantRNE_48U_24U_else_and_tmp;
  wire IsNaN_8U_23U_1_nor_3_tmp;
  wire IsNaN_8U_23U_1_nor_2_tmp;
  wire IsNaN_8U_23U_1_nor_1_tmp;
  wire IsNaN_8U_23U_1_nor_tmp;
  wire or_tmp_1;
  wire not_tmp_2;
  wire or_tmp_12;
  wire or_tmp_15;
  wire not_tmp_8;
  wire or_tmp_26;
  wire or_tmp_29;
  wire not_tmp_12;
  wire or_tmp_40;
  wire not_tmp_15;
  wire or_tmp_46;
  wire or_tmp_51;
  wire or_tmp_59;
  wire or_tmp_75;
  wire or_tmp_91;
  wire or_tmp_107;
  wire or_tmp_123;
  wire or_tmp_128;
  wire or_tmp_132;
  wire or_tmp_133;
  wire or_tmp_146;
  wire or_tmp_167;
  wire or_tmp_173;
  wire mux_tmp_46;
  wire mux_tmp_48;
  wire not_tmp_54;
  wire not_tmp_55;
  wire or_tmp_211;
  wire or_tmp_216;
  wire or_tmp_235;
  wire or_tmp_252;
  wire or_tmp_256;
  wire mux_tmp_78;
  wire not_tmp_81;
  wire not_tmp_82;
  wire or_tmp_291;
  wire or_tmp_296;
  wire or_tmp_315;
  wire or_tmp_332;
  wire or_tmp_336;
  wire mux_tmp_109;
  wire not_tmp_106;
  wire not_tmp_107;
  wire or_tmp_371;
  wire or_tmp_376;
  wire not_tmp_121;
  wire or_tmp_395;
  wire or_tmp_411;
  wire or_tmp_415;
  wire mux_tmp_140;
  wire not_tmp_129;
  wire not_tmp_130;
  wire or_tmp_461;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_11;
  wire and_dcpl_14;
  wire or_tmp_517;
  wire and_tmp_5;
  wire and_dcpl_22;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire or_dcpl_8;
  wire and_dcpl_30;
  wire or_dcpl_13;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_37;
  wire or_dcpl_40;
  wire or_dcpl_50;
  wire or_dcpl_53;
  wire or_dcpl_63;
  wire or_dcpl_66;
  wire or_dcpl_75;
  wire or_dcpl_81;
  wire or_dcpl_87;
  wire or_dcpl_93;
  wire or_dcpl_96;
  wire or_dcpl_99;
  wire or_dcpl_102;
  wire or_dcpl_105;
  wire or_dcpl_108;
  wire or_dcpl_110;
  wire or_dcpl_125;
  wire or_tmp_587;
  wire or_tmp_588;
  wire or_tmp_591;
  reg IsZero_8U_23U_land_1_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm_5;
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_1_sva;
  reg [7:0] FpMul_8U_23U_p_expo_1_sva_1;
  reg FpMantRNE_48U_24U_else_carry_1_sva;
  reg IsZero_8U_23U_land_2_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm_5;
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_2_sva;
  reg [7:0] FpMul_8U_23U_p_expo_2_sva_1;
  reg FpMantRNE_48U_24U_else_carry_2_sva;
  reg IsZero_8U_23U_land_3_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm_5;
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_3_sva;
  reg [7:0] FpMul_8U_23U_p_expo_3_sva_1;
  reg FpMantRNE_48U_24U_else_carry_3_sva;
  reg IsZero_8U_23U_land_lpi_1_dfm;
  reg IsZero_8U_23U_1_land_lpi_1_dfm_5;
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  reg [47:0] FpMul_8U_23U_p_mant_p1_sva;
  reg [7:0] FpMul_8U_23U_p_expo_sva_1;
  reg FpMantRNE_48U_24U_else_carry_sva;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg mul_mul_land_1_lpi_1_dfm_2;
  reg mul_mul_land_1_lpi_1_dfm_5;
  reg mul_mul_land_1_lpi_1_dfm_6;
  reg mul_mul_land_2_lpi_1_dfm_2;
  reg mul_mul_land_2_lpi_1_dfm_5;
  reg mul_mul_land_2_lpi_1_dfm_6;
  reg mul_mul_land_3_lpi_1_dfm_2;
  reg mul_mul_land_3_lpi_1_dfm_5;
  reg mul_mul_land_3_lpi_1_dfm_6;
  reg mul_mul_land_lpi_1_dfm_2;
  reg mul_mul_land_lpi_1_dfm_5;
  reg mul_mul_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  reg cfg_mul_src_1_sva_1;
  reg [31:0] cfg_mul_op_1_sva_1;
  reg [9:0] cfg_truncate_1_sva_1;
  reg [9:0] cfg_truncate_1_sva_3;
  reg [127:0] MulIn_data_sva_1;
  reg [127:0] MulIn_data_sva_132;
  reg [127:0] MulIn_data_sva_133;
  reg io_read_cfg_mul_bypass_rsc_svs_5;
  reg IsZero_8U_23U_land_1_lpi_1_dfm_4;
  reg IsZero_8U_23U_land_1_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg [7:0] FpMul_8U_23U_p_expo_1_sva_5;
  reg FpMantRNE_48U_24U_else_carry_1_sva_2;
  reg mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsZero_8U_23U_land_2_lpi_1_dfm_4;
  reg IsZero_8U_23U_land_2_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg [7:0] FpMul_8U_23U_p_expo_2_sva_5;
  reg FpMantRNE_48U_24U_else_carry_2_sva_2;
  reg mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsZero_8U_23U_land_3_lpi_1_dfm_4;
  reg IsZero_8U_23U_land_3_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg [7:0] FpMul_8U_23U_p_expo_3_sva_5;
  reg FpMantRNE_48U_24U_else_carry_3_sva_2;
  reg mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  reg IsZero_8U_23U_land_lpi_1_dfm_4;
  reg IsZero_8U_23U_land_lpi_1_dfm_6;
  reg IsZero_8U_23U_1_land_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  reg [7:0] FpMul_8U_23U_p_expo_sva_5;
  reg FpMantRNE_48U_24U_else_carry_sva_2;
  reg mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  reg cfg_mul_src_1_sva_st;
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st;
  reg mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  reg [22:0] mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  reg mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st;
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2;
  reg [63:0] mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm;
  reg [63:0] mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2;
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st;
  reg mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_12_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2;
  reg [22:0] mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  reg mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st;
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2;
  reg [63:0] mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm;
  reg [63:0] mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2;
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st;
  reg mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_13_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2;
  reg [22:0] mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  reg mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st;
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2;
  reg [63:0] mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm;
  reg [63:0] mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2;
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  reg mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm;
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2;
  reg FpMul_8U_23U_FpMul_8U_23U_and_14_itm;
  reg FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2;
  reg [22:0] mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  reg mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st;
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm;
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2;
  reg [63:0] mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm;
  reg [63:0] mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2;
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  reg FpMul_8U_23U_mux_49_itm_3;
  reg FpMul_8U_23U_mux_49_itm_4;
  reg FpMul_8U_23U_mux_36_itm_3;
  reg FpMul_8U_23U_mux_36_itm_4;
  reg FpMul_8U_23U_mux_23_itm_3;
  reg FpMul_8U_23U_mux_23_itm_4;
  reg FpMul_8U_23U_mux_10_itm_3;
  reg FpMul_8U_23U_mux_10_itm_4;
  reg io_read_cfg_mul_bypass_rsc_svs_st_1;
  reg cfg_mul_src_1_sva_st_1;
  reg mul_mul_land_1_lpi_1_dfm_st_1;
  reg io_read_cfg_mul_bypass_rsc_svs_st_4;
  reg mul_mul_land_1_lpi_1_dfm_st_4;
  reg mul_mul_land_1_lpi_1_dfm_st_5;
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st_4;
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3;
  reg mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_1;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  reg mul_mul_land_2_lpi_1_dfm_st_1;
  reg mul_mul_land_2_lpi_1_dfm_st_4;
  reg mul_mul_land_2_lpi_1_dfm_st_5;
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st_4;
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3;
  reg mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_1;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  reg mul_mul_land_3_lpi_1_dfm_st_1;
  reg mul_mul_land_3_lpi_1_dfm_st_4;
  reg mul_mul_land_3_lpi_1_dfm_st_5;
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st_4;
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3;
  reg mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_1;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  reg mul_mul_land_lpi_1_dfm_st_1;
  reg mul_mul_land_lpi_1_dfm_st_4;
  reg mul_mul_land_lpi_1_dfm_st_5;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  reg mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3;
  reg mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_1;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  reg [30:0] else_MulOp_data_0_lpi_1_dfm_2_30_0_1;
  reg [30:0] else_MulOp_data_1_lpi_1_dfm_2_30_0_1;
  reg [30:0] else_MulOp_data_2_lpi_1_dfm_2_30_0_1;
  reg [30:0] else_MulOp_data_3_lpi_1_dfm_2_30_0_1;
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1;
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1;
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1;
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1;
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1;
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1;
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1;
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1;
  wire [7:0] else_mux_3_tmp_30_23;
  wire [7:0] else_mux_2_tmp_30_23;
  wire [7:0] else_mux_1_tmp_30_23;
  wire [7:0] else_mux_tmp_30_23;
  wire mul_mul_else_unequal_tmp_1;
  wire FpMul_8U_23U_is_inf_1_lpi_1_dfm_2;
  wire [7:0] FpMul_8U_23U_o_expo_lpi_1_dfm;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  wire [7:0] FpMul_8U_23U_o_expo_3_lpi_1_dfm;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  wire [7:0] FpMul_8U_23U_o_expo_2_lpi_1_dfm;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  wire [7:0] FpMul_8U_23U_o_expo_1_lpi_1_dfm;
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp;
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva;
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva;
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva;
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva;
  wire [47:0] FpMul_8U_23U_p_mant_p1_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_3_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_2_sva_mx1;
  wire [47:0] FpMul_8U_23U_p_mant_p1_1_sva_mx1;
  wire [30:0] else_MulOp_data_3_lpi_1_dfm_mx0_30_0;
  wire [30:0] else_MulOp_data_2_lpi_1_dfm_mx0_30_0;
  wire [30:0] else_MulOp_data_1_lpi_1_dfm_mx0_30_0;
  wire [30:0] else_MulOp_data_0_lpi_1_dfm_mx0_30_0;
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva;
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva;
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva;
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva;
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva;
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva;
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva;
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva;
  wire and_142_m1c;
  wire and_140_m1c;
  wire and_138_m1c;
  wire and_136_m1c;
  wire mul_mul_and_21_m1c;
  wire mul_mul_and_19_m1c;
  wire mul_mul_and_17_m1c;
  wire mul_mul_and_m1c;
  wire chn_mul_out_and_1_cse;
  wire chn_mul_out_and_cse;
  reg reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse;
  wire or_27_cse;
  wire or_74_cse;
  wire nor_20_cse;
  wire nor_301_cse;
  wire nor_277_cse;
  wire nor_31_cse;
  wire nor_282_cse;
  wire nor_264_cse;
  wire nor_267_cse;
  wire nor_241_cse;
  wire nor_49_cse;
  wire nor_245_cse;
  wire nor_227_cse;
  wire nor_230_cse;
  wire nor_204_cse;
  wire nor_68_cse;
  wire nor_208_cse;
  wire nor_190_cse;
  wire nor_193_cse;
  wire nor_170_cse;
  wire nor_86_cse;
  wire nor_174_cse;
  reg reg_chn_mul_out_rsci_ld_core_psct_cse;
  wire IsNaN_8U_23U_aelse_and_cse;
  wire MulIn_data_and_cse;
  wire FpMul_8U_23U_p_expo_and_cse;
  wire else_MulOp_data_and_1_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_cse;
  wire nor_143_cse;
  wire FpMul_8U_23U_p_expo_and_1_cse;
  wire else_MulOp_data_and_3_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse;
  wire FpMul_8U_23U_p_expo_and_2_cse;
  wire else_MulOp_data_and_5_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse;
  wire or_430_cse;
  wire FpMul_8U_23U_p_expo_and_3_cse;
  wire else_MulOp_data_and_7_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse;
  wire or_468_cse;
  wire IsNaN_8U_23U_aelse_and_4_cse;
  wire IsNaN_8U_23U_aelse_and_5_cse;
  wire IsNaN_8U_23U_aelse_and_6_cse;
  wire IsNaN_8U_23U_aelse_and_7_cse;
  wire or_469_cse;
  wire or_482_cse;
  wire or_490_cse;
  wire nand_48_cse;
  wire nand_45_cse;
  wire nand_42_cse;
  wire nor_118_cse;
  wire nor_117_cse;
  wire nor_116_cse;
  wire nor_115_cse;
  wire or_189_cse;
  wire nor_348_cse;
  wire nor_347_cse;
  wire nor_346_cse;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0;
  wire [45:0] FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0;
  wire and_135_rgt;
  wire mul_mul_if_and_6_rgt;
  wire mul_mul_if_and_7_rgt;
  wire and_137_rgt;
  wire mul_mul_if_and_4_rgt;
  wire mul_mul_if_and_5_rgt;
  wire and_139_rgt;
  wire mul_mul_if_and_2_rgt;
  wire mul_mul_if_and_3_rgt;
  wire and_141_rgt;
  wire mul_mul_if_and_rgt;
  wire mul_mul_if_and_1_rgt;
  wire and_146_rgt;
  wire and_150_rgt;
  wire and_154_rgt;
  wire and_158_rgt;
  wire mux_7_itm;
  wire mux_12_itm;
  wire mux_17_itm;
  wire mux_22_itm;
  wire mux_94_itm;
  wire mux_125_itm;
  wire chn_mul_in_rsci_ld_core_psct_mx0c0;
  wire chn_mul_op_rsci_ld_core_psct_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire [7:0] FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_1_sva_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0;
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_2_sva_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0;
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_3_sva_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0;
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  wire [7:0] FpMul_8U_23U_p_expo_sva_1_mx0w0;
  wire [8:0] nl_FpMul_8U_23U_p_expo_sva_1_mx0w0;
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0;
  wire FpMantRNE_48U_24U_else_carry_sva_mx0w0;
  wire FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0;
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  wire main_stage_v_1_mx0c1;
  wire IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0;
  wire IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0;
  wire IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0;
  wire IsZero_8U_23U_land_lpi_1_dfm_mx1w0;
  wire mul_mul_land_lpi_1_dfm_mx1w0;
  wire mul_mul_land_3_lpi_1_dfm_mx1w0;
  wire mul_mul_land_2_lpi_1_dfm_mx1w0;
  wire mul_mul_land_1_lpi_1_dfm_mx1w0;
  wire cfg_mul_src_1_sva_st_1_mx0c1;
  wire FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
  wire FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0;
  wire [63:0] mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  wire [63:0] mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  wire [63:0] mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  wire [63:0] mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  wire IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
  wire [22:0] FpMul_8U_23U_o_mant_1_lpi_1_dfm_3;
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva;
  wire [22:0] FpMul_8U_23U_o_mant_2_lpi_1_dfm_3;
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva;
  wire [22:0] FpMul_8U_23U_o_mant_3_lpi_1_dfm_3;
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva;
  wire [22:0] FpMul_8U_23U_o_mant_lpi_1_dfm_3;
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva;
  wire mul_mul_mul_mul_nor_6_m1c;
  wire mul_mul_mul_mul_nor_4_m1c;
  wire mul_mul_mul_mul_nor_2_m1c;
  wire mul_mul_mul_mul_nor_m1c;
  wire [7:0] FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0;
  wire FpMul_8U_23U_lor_9_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0;
  wire FpMul_8U_23U_lor_10_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0;
  wire FpMul_8U_23U_lor_11_lpi_1_dfm;
  wire [7:0] FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0;
  wire FpMul_8U_23U_lor_2_lpi_1_dfm;
  wire [31:0] else_MulOp_data_0_lpi_1_dfm_mx1;
  wire [31:0] else_MulOp_data_1_lpi_1_dfm_mx1;
  wire [31:0] else_MulOp_data_2_lpi_1_dfm_mx1;
  wire [31:0] else_MulOp_data_3_lpi_1_dfm_mx1;
  wire or_11_cse;
  wire or_12_cse;
  wire or_13_cse;
  wire or_14_cse;
  wire or_15_cse;
  wire or_16_cse;
  wire asn_156;
  wire asn_158;
  wire asn_160;
  wire asn_162;
  wire asn_164;
  wire asn_166;
  wire asn_168;
  wire asn_170;
  wire IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse;
  wire else_MulOp_data_and_8_cse;
  wire else_MulOp_data_and_9_cse;
  wire else_MulOp_data_and_10_cse;
  wire else_MulOp_data_and_11_cse;
  wire mul_mul_aelse_and_cse;
  wire MulIn_data_and_1_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse;
  wire FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse;
  wire MulIn_data_and_2_cse;
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
  wire IsNaN_8U_23U_aelse_and_17_cse;
  wire IsNaN_8U_23U_1_aelse_and_cse;
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
  wire IsNaN_8U_23U_aelse_and_19_cse;
  wire IsNaN_8U_23U_1_aelse_and_1_cse;
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
  wire IsNaN_8U_23U_aelse_and_21_cse;
  wire IsNaN_8U_23U_1_aelse_and_2_cse;
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse;
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
  wire IsNaN_8U_23U_aelse_and_23_cse;
  wire IsNaN_8U_23U_1_aelse_and_3_cse;
  wire mul_mul_aelse_and_12_cse;
  wire IsNaN_8U_23U_aelse_and_24_cse;
  wire IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse;
  wire mul_mul_aelse_and_19_cse;
  wire FpMantRNE_48U_24U_else_and_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse;
  wire FpMantRNE_48U_24U_else_and_9_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse;
  wire FpMantRNE_48U_24U_else_and_11_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse;
  wire FpMantRNE_48U_24U_else_and_13_cse;
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse;
  wire IsNaN_8U_23U_aelse_and_25_cse;
  wire IsNaN_8U_23U_aelse_and_26_cse;
  wire IsNaN_8U_23U_aelse_and_27_cse;
  wire FpMul_8U_23U_oelse_1_and_4_cse;
  wire FpMul_8U_23U_oelse_1_and_5_cse;
  wire FpMul_8U_23U_oelse_1_and_6_cse;
  wire FpMul_8U_23U_oelse_1_and_7_cse;
  wire mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  wire mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  wire mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  wire mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  wire mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  wire mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;

  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] and_59;
  wire[0:0] oWidth_aWidth_bWidth_prb;
  wire[0:0] and_61;
  wire[0:0] iMantWidth_oMantWidth_prb_1;
  wire[0:0] and_63;
  wire[0:0] oWidth_aWidth_bWidth_prb_1;
  wire[0:0] and_65;
  wire[0:0] iMantWidth_oMantWidth_prb_2;
  wire[0:0] and_67;
  wire[0:0] oWidth_aWidth_bWidth_prb_2;
  wire[0:0] and_69;
  wire[0:0] iMantWidth_oMantWidth_prb_3;
  wire[0:0] and_71;
  wire[0:0] oWidth_aWidth_bWidth_prb_3;
  wire[0:0] and_73;
  wire[0:0] mul_mul_mux_108_nl;
  wire[0:0] mul_mul_else_mux_26_nl;
  wire[0:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  wire[21:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  wire[21:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] nor_3_nl;
  wire[7:0] FpMul_8U_23U_FpMul_8U_23U_and_15_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_4_nl;
  wire[7:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  wire[7:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  wire[0:0] and_358_nl;
  wire[0:0] and_359_nl;
  wire[0:0] or_839_nl;
  wire[0:0] mul_mul_mux_109_nl;
  wire[0:0] mul_mul_else_mux_23_nl;
  wire[0:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] mul_mul_mux_110_nl;
  wire[0:0] mul_mul_else_mux_53_nl;
  wire[0:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  wire[21:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  wire[21:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] nor_2_nl;
  wire[7:0] FpMul_8U_23U_FpMul_8U_23U_and_16_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_5_nl;
  wire[7:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  wire[7:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  wire[0:0] and_356_nl;
  wire[0:0] and_357_nl;
  wire[0:0] or_838_nl;
  wire[0:0] mul_mul_mux_111_nl;
  wire[0:0] mul_mul_else_mux_50_nl;
  wire[0:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] mul_mul_mux_112_nl;
  wire[0:0] mul_mul_else_mux_80_nl;
  wire[0:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  wire[21:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  wire[21:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] nor_1_nl;
  wire[7:0] FpMul_8U_23U_FpMul_8U_23U_and_17_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_6_nl;
  wire[7:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  wire[7:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  wire[0:0] and_354_nl;
  wire[0:0] and_355_nl;
  wire[0:0] or_837_nl;
  wire[0:0] mul_mul_mux_113_nl;
  wire[0:0] mul_mul_else_mux_77_nl;
  wire[0:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] mul_mul_mux_114_nl;
  wire[0:0] mul_mul_else_mux_107_nl;
  wire[0:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  wire[21:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  wire[21:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] nor_6_nl;
  wire[7:0] FpMul_8U_23U_FpMul_8U_23U_and_18_nl;
  wire[0:0] FpMul_8U_23U_oelse_2_not_7_nl;
  wire[7:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  wire[7:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  wire[0:0] and_352_nl;
  wire[0:0] and_353_nl;
  wire[0:0] or_836_nl;
  wire[0:0] mul_mul_mux_115_nl;
  wire[0:0] mul_mul_else_mux_104_nl;
  wire[0:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_28_nl;
  wire[0:0] or_31_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] or_42_nl;
  wire[0:0] or_45_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] or_56_nl;
  wire[0:0] or_59_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] or_67_nl;
  wire[0:0] or_70_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] nor_319_nl;
  wire[0:0] nor_320_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] nor_315_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] nor_311_nl;
  wire[0:0] nor_312_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] and_344_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] or_142_nl;
  wire[0:0] or_143_nl;
  wire[0:0] or_831_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] or_147_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] mux_41_nl;
  wire[0:0] or_153_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] nor_297_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] or_165_nl;
  wire[0:0] or_166_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] or_169_nl;
  wire[0:0] nor_294_nl;
  wire[0:0] mux_50_nl;
  wire[0:0] nor_290_nl;
  wire[0:0] nor_291_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] or_181_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] or_185_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] or_211_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] nor_276_nl;
  wire[0:0] nor_278_nl;
  wire[0:0] or_210_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] and_343_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] nor_269_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] nor_272_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] nor_263_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] or_227_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] or_230_nl;
  wire[0:0] or_231_nl;
  wire[0:0] or_830_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] or_235_nl;
  wire[0:0] nor_266_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] nor_268_nl;
  wire[0:0] and_342_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] nor_260_nl;
  wire[0:0] nor_261_nl;
  wire[0:0] nor_262_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] or_254_nl;
  wire[0:0] or_255_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] or_258_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] nor_253_nl;
  wire[0:0] nor_254_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] or_270_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] and_340_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] nor_238_nl;
  wire[0:0] nor_239_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] nor_240_nl;
  wire[0:0] nor_242_nl;
  wire[0:0] or_292_nl;
  wire[0:0] nor_243_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] and_339_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] nor_232_nl;
  wire[0:0] nor_234_nl;
  wire[0:0] nor_235_nl;
  wire[0:0] nor_236_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] nor_226_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] or_307_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] or_310_nl;
  wire[0:0] or_311_nl;
  wire[0:0] or_829_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] or_315_nl;
  wire[0:0] nor_229_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] nor_231_nl;
  wire[0:0] and_338_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] nor_223_nl;
  wire[0:0] nor_224_nl;
  wire[0:0] nor_225_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] nor_218_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] or_334_nl;
  wire[0:0] or_335_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] or_338_nl;
  wire[0:0] nor_220_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] nor_216_nl;
  wire[0:0] nor_217_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] or_350_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] and_336_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_201_nl;
  wire[0:0] nor_202_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] nand_29_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] nor_203_nl;
  wire[0:0] nor_205_nl;
  wire[0:0] or_372_nl;
  wire[0:0] nor_206_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] and_335_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] nor_195_nl;
  wire[0:0] nor_197_nl;
  wire[0:0] nor_198_nl;
  wire[0:0] nor_199_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] nor_189_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] or_387_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] or_390_nl;
  wire[0:0] or_391_nl;
  wire[0:0] or_828_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] or_395_nl;
  wire[0:0] nor_192_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] nor_194_nl;
  wire[0:0] and_334_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] nor_186_nl;
  wire[0:0] nor_187_nl;
  wire[0:0] nor_188_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] nor_181_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] or_414_nl;
  wire[0:0] or_415_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] or_418_nl;
  wire[0:0] nor_183_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] or_429_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] or_424_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] or_436_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] and_332_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] nor_167_nl;
  wire[0:0] nor_168_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] nor_169_nl;
  wire[0:0] nor_171_nl;
  wire[0:0] or_453_nl;
  wire[0:0] nor_172_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] and_331_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] nor_161_nl;
  wire[0:0] nor_163_nl;
  wire[0:0] nor_164_nl;
  wire[0:0] nor_165_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] or_467_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] or_480_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] or_488_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] or_496_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] or_511_nl;
  wire[0:0] nor_144_nl;
  wire[0:0] or_509_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] and_39_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] or_515_nl;
  wire[0:0] nor_100_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] or_519_nl;
  wire[0:0] nor_142_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] and_40_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] or_523_nl;
  wire[0:0] nor_102_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] or_527_nl;
  wire[0:0] nor_140_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] and_41_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] or_531_nl;
  wire[0:0] nor_104_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] or_535_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] nor_107_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] and_328_nl;
  wire[0:0] FpMul_8U_23U_oelse_1_mux_20_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] nor_136_nl;
  wire[0:0] nor_137_nl;
  wire[0:0] or_540_nl;
  wire[0:0] nor_138_nl;
  wire[0:0] mul_mul_1_FpMul_8U_23U_xor_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] nor_134_nl;
  wire[0:0] nor_135_nl;
  wire[0:0] FpMul_8U_23U_oelse_1_mux_21_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] nor_131_nl;
  wire[0:0] nor_132_nl;
  wire[0:0] or_551_nl;
  wire[0:0] nor_133_nl;
  wire[0:0] mul_mul_2_FpMul_8U_23U_xor_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] nor_129_nl;
  wire[0:0] nor_130_nl;
  wire[0:0] FpMul_8U_23U_oelse_1_mux_22_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] nor_126_nl;
  wire[0:0] nor_127_nl;
  wire[0:0] or_561_nl;
  wire[0:0] nor_128_nl;
  wire[0:0] mul_mul_3_FpMul_8U_23U_xor_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] nor_124_nl;
  wire[0:0] nor_125_nl;
  wire[0:0] FpMul_8U_23U_oelse_1_mux_23_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] nor_121_nl;
  wire[0:0] nor_122_nl;
  wire[0:0] or_571_nl;
  wire[0:0] nor_123_nl;
  wire[0:0] mul_mul_4_FpMul_8U_23U_xor_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] nor_119_nl;
  wire[0:0] nor_120_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] nor_159_nl;
  wire[0:0] or_473_nl;
  wire[0:0] or_474_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] nor_157_nl;
  wire[0:0] or_486_nl;
  wire[0:0] or_487_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] nor_155_nl;
  wire[0:0] or_494_nl;
  wire[0:0] or_495_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] or_498_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] nor_153_nl;
  wire[0:0] or_502_nl;
  wire[0:0] or_503_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_2_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_2_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_3_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_3_nl;
  wire[7:0] FpMul_8U_23U_else_2_else_acc_4_nl;
  wire[8:0] nl_FpMul_8U_23U_else_2_else_acc_4_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_7_nl;
  wire[8:0] mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_6_nl;
  wire[8:0] mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_5_nl;
  wire[8:0] mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  wire[0:0] FpMul_8U_23U_p_mant_p1_and_4_nl;
  wire[8:0] mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  wire[9:0] nl_mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  wire[8:0] mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  wire[9:0] nl_mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  wire[22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_4_nl;
  wire[22:0] FpMul_8U_23U_nor_nl;
  wire[22:0] mux_237_nl;
  wire[22:0] mul_mul_1_FpMantRNE_48U_24U_else_acc_nl;
  wire[23:0] nl_mul_mul_1_FpMantRNE_48U_24U_else_acc_nl;
  wire[0:0] or_nl;
  wire[0:0] FpMul_8U_23U_FpMul_8U_23U_nor_nl;
  wire[0:0] FpMul_8U_23U_and_1_nl;
  wire[22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_5_nl;
  wire[22:0] FpMul_8U_23U_nor_4_nl;
  wire[22:0] mux_238_nl;
  wire[22:0] mul_mul_2_FpMantRNE_48U_24U_else_acc_nl;
  wire[23:0] nl_mul_mul_2_FpMantRNE_48U_24U_else_acc_nl;
  wire[0:0] or_840_nl;
  wire[0:0] FpMul_8U_23U_FpMul_8U_23U_nor_1_nl;
  wire[0:0] FpMul_8U_23U_and_3_nl;
  wire[22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_6_nl;
  wire[22:0] FpMul_8U_23U_nor_5_nl;
  wire[22:0] mux_239_nl;
  wire[22:0] mul_mul_3_FpMantRNE_48U_24U_else_acc_nl;
  wire[23:0] nl_mul_mul_3_FpMantRNE_48U_24U_else_acc_nl;
  wire[0:0] or_841_nl;
  wire[0:0] FpMul_8U_23U_FpMul_8U_23U_nor_2_nl;
  wire[0:0] FpMul_8U_23U_and_5_nl;
  wire[22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_7_nl;
  wire[22:0] FpMul_8U_23U_nor_6_nl;
  wire[22:0] mux_240_nl;
  wire[22:0] mul_mul_4_FpMantRNE_48U_24U_else_acc_nl;
  wire[23:0] nl_mul_mul_4_FpMantRNE_48U_24U_else_acc_nl;
  wire[0:0] or_842_nl;
  wire[0:0] FpMul_8U_23U_FpMul_8U_23U_nor_3_nl;
  wire[0:0] FpMul_8U_23U_and_7_nl;
  wire[7:0] mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_8U_23U_FpMul_8U_23U_nor_4_nl;
  wire[0:0] FpMul_8U_23U_or_4_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl;
  wire[7:0] mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_8U_23U_or_5_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl;
  wire[7:0] mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_8U_23U_or_6_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl;
  wire[7:0] mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[8:0] nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_8U_23U_or_7_nl;
  wire[0:0] FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl;
  wire[9:0] mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_nl;
  wire[9:0] mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_1_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_1_nl;
  wire[9:0] mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_2_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_2_nl;
  wire[9:0] mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  wire[10:0] nl_mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  wire[8:0] FpMul_8U_23U_oelse_1_acc_3_nl;
  wire[9:0] nl_FpMul_8U_23U_oelse_1_acc_3_nl;
  wire[0:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  wire[0:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  wire[0:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  wire[0:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  wire[7:0] mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] or_743_nl;
  wire[7:0] mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] or_744_nl;
  wire[7:0] mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] or_745_nl;
  wire[7:0] mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[8:0] nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] or_19_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] or_26_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] or_34_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] or_40_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] or_48_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] or_54_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_321_nl;
  wire[0:0] nor_322_nl;
  wire[0:0] nor_323_nl;
  wire[0:0] or_65_nl;
  wire[0:0] or_187_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] nor_288_nl;
  wire[0:0] nor_289_nl;
  wire[0:0] or_193_nl;
  wire[0:0] nor_283_nl;
  wire[0:0] nor_284_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] nor_251_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] nor_246_nl;
  wire[0:0] nor_247_nl;
  wire[0:0] nor_211_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] nor_212_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] nor_214_nl;
  wire[0:0] nor_215_nl;
  wire[0:0] nor_209_nl;
  wire[0:0] nor_210_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] or_435_nl;
  wire[0:0] nor_177_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] nor_179_nl;
  wire[0:0] nor_180_nl;
  wire[0:0] nor_175_nl;
  wire[0:0] nor_176_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [1086:0] nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  assign nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = {mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2
      , {512'b0 , 511'b0}};
  wire [9:0] nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  assign nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  wire [1086:0] nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  assign nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = {mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2
      , {512'b0 , 511'b0}};
  wire [9:0] nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  assign nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  wire [1086:0] nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  assign nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = {mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2
      , {512'b0 , 511'b0}};
  wire [9:0] nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  assign nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  wire [1086:0] nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  assign nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = {mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2
      , {512'b0 , 511'b0}};
  wire [9:0] nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  assign nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  wire [127:0] nl_Y_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d;
  assign nl_Y_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d = {chn_mul_out_rsci_d_127
      , chn_mul_out_rsci_d_126_119 , chn_mul_out_rsci_d_118_97 , chn_mul_out_rsci_d_96
      , chn_mul_out_rsci_d_95 , chn_mul_out_rsci_d_94_87 , chn_mul_out_rsci_d_86_65
      , chn_mul_out_rsci_d_64 , chn_mul_out_rsci_d_63 , chn_mul_out_rsci_d_62_55
      , chn_mul_out_rsci_d_54_33 , chn_mul_out_rsci_d_32 , chn_mul_out_rsci_d_31
      , chn_mul_out_rsci_d_30_23 , chn_mul_out_rsci_d_22_1 , chn_mul_out_rsci_d_0};
  SDP_Y_CORE_mgc_shift_r_v4 #(.width_a(32'sd1087),
  .signd_a(32'sd1),
  .width_s(32'sd10),
  .width_z(32'sd1087)) mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a[1086:0]),
      .s(nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s[9:0]),
      .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva)
    );
  SDP_Y_CORE_mgc_shift_r_v4 #(.width_a(32'sd1087),
  .signd_a(32'sd1),
  .width_s(32'sd10),
  .width_z(32'sd1087)) mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a[1086:0]),
      .s(nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s[9:0]),
      .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva)
    );
  SDP_Y_CORE_mgc_shift_r_v4 #(.width_a(32'sd1087),
  .signd_a(32'sd1),
  .width_s(32'sd10),
  .width_z(32'sd1087)) mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a[1086:0]),
      .s(nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s[9:0]),
      .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva)
    );
  SDP_Y_CORE_mgc_shift_r_v4 #(.width_a(32'sd1087),
  .signd_a(32'sd1),
  .width_s(32'sd10),
  .width_z(32'sd1087)) mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a[1086:0]),
      .s(nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s[9:0]),
      .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci Y_mul_core_chn_mul_in_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsc_z(chn_mul_in_rsc_z),
      .chn_mul_in_rsc_vz(chn_mul_in_rsc_vz),
      .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_mul_in_rsci_iswt0(chn_mul_in_rsci_iswt0),
      .chn_mul_in_rsci_bawt(chn_mul_in_rsci_bawt),
      .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
      .chn_mul_in_rsci_ld_core_psct(chn_mul_in_rsci_ld_core_psct),
      .chn_mul_in_rsci_d_mxwt(chn_mul_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci Y_mul_core_chn_mul_op_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
      .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
      .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_op_rsci_iswt0(chn_mul_op_rsci_iswt0),
      .chn_mul_op_rsci_bawt(chn_mul_op_rsci_bawt),
      .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
      .chn_mul_op_rsci_ld_core_psct(chn_mul_op_rsci_ld_core_psct),
      .chn_mul_op_rsci_d_mxwt(chn_mul_op_rsci_d_mxwt)
    );
  SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci Y_mul_core_chn_mul_out_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_out_rsc_z(chn_mul_out_rsc_z),
      .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz),
      .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_mul_out_rsci_iswt0(chn_mul_out_rsci_iswt0),
      .chn_mul_out_rsci_bawt(chn_mul_out_rsci_bawt),
      .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp),
      .chn_mul_out_rsci_ld_core_psct(reg_chn_mul_out_rsci_ld_core_psct_cse),
      .chn_mul_out_rsci_d(nl_Y_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d[127:0])
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz),
      .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_bypass_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_bypass_rsc_triosy_obj_bawt(cfg_mul_bypass_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz),
      .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_prelu_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_prelu_rsc_triosy_obj_bawt(cfg_mul_prelu_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj Y_mul_core_cfg_mul_src_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz),
      .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_src_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_src_rsc_triosy_obj_bawt(cfg_mul_src_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj Y_mul_core_cfg_mul_op_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz),
      .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_mul_op_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_mul_op_rsc_triosy_obj_bawt(cfg_mul_op_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj Y_mul_core_cfg_truncate_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_truncate_rsc_triosy_lz(cfg_truncate_rsc_triosy_lz),
      .cfg_truncate_rsc_triosy_obj_oswt(cfg_truncate_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_truncate_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_truncate_rsc_triosy_obj_bawt(cfg_truncate_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_mul_core_staller Y_mul_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
      .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp)
    );
  SDP_Y_CORE_Y_mul_core_core_fsm Y_mul_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_59 = and_dcpl_4 & and_dcpl_3 & (fsm_output[1]);
  assign iMantWidth_oMantWidth_prb = MUX1HOT_s_1_1_2(1'b1, and_59);
  // assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
  // PSL mul_mul_1_Y_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign and_61 = and_dcpl_4 & and_dcpl_6 & (fsm_output[1]);
  assign oWidth_aWidth_bWidth_prb = MUX1HOT_s_1_1_2(1'b1, and_61);
  // assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
  // PSL mul_mul_1_Y_mul_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth : assert { oWidth_aWidth_bWidth_prb } @rose(nvdla_core_clk);
  assign and_63 = and_dcpl_8 & and_dcpl_3 & (fsm_output[1]);
  assign iMantWidth_oMantWidth_prb_1 = MUX1HOT_s_1_1_2(1'b1, and_63);
  // assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
  // PSL mul_mul_2_Y_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_1 } @rose(nvdla_core_clk);
  assign and_65 = and_dcpl_8 & and_dcpl_6 & (fsm_output[1]);
  assign oWidth_aWidth_bWidth_prb_1 = MUX1HOT_s_1_1_2(1'b1, and_65);
  // assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
  // PSL mul_mul_2_Y_mul_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth : assert { oWidth_aWidth_bWidth_prb_1 } @rose(nvdla_core_clk);
  assign and_67 = and_dcpl_11 & and_dcpl_3 & (fsm_output[1]);
  assign iMantWidth_oMantWidth_prb_2 = MUX1HOT_s_1_1_2(1'b1, and_67);
  // assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
  // PSL mul_mul_3_Y_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_2 } @rose(nvdla_core_clk);
  assign and_69 = and_dcpl_11 & and_dcpl_6 & (fsm_output[1]);
  assign oWidth_aWidth_bWidth_prb_2 = MUX1HOT_s_1_1_2(1'b1, and_69);
  // assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
  // PSL mul_mul_3_Y_mul_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth : assert { oWidth_aWidth_bWidth_prb_2 } @rose(nvdla_core_clk);
  assign and_71 = and_dcpl_14 & and_dcpl_3 & (fsm_output[1]);
  assign iMantWidth_oMantWidth_prb_3 = MUX1HOT_s_1_1_2(1'b1, and_71);
  // assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
  // PSL mul_mul_4_Y_mul_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_3 } @rose(nvdla_core_clk);
  assign and_73 = and_dcpl_14 & and_dcpl_6 & (fsm_output[1]);
  assign oWidth_aWidth_bWidth_prb_3 = MUX1HOT_s_1_1_2(1'b1, and_73);
  // assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
  // PSL mul_mul_4_Y_mul_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth : assert { oWidth_aWidth_bWidth_prb_3 } @rose(nvdla_core_clk);
  assign chn_mul_out_and_cse = core_wen & ((main_stage_v_3 & io_read_cfg_mul_bypass_rsc_svs_5
      & or_74_cse) | and_dcpl_22);
  assign chn_mul_out_and_1_cse = core_wen & (~(and_dcpl_23 | (~ main_stage_v_3)));
  assign mul_mul_and_m1c = (~ IsNaN_8U_23U_land_1_lpi_1_dfm_8) & mul_mul_mul_mul_nor_m1c
      & (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign mul_mul_and_17_m1c = (~ IsNaN_8U_23U_land_2_lpi_1_dfm_8) & mul_mul_mul_mul_nor_2_m1c
      & (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign mul_mul_and_19_m1c = (~ IsNaN_8U_23U_land_3_lpi_1_dfm_8) & mul_mul_mul_mul_nor_4_m1c
      & (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign mul_mul_and_21_m1c = (~ IsNaN_8U_23U_land_lpi_1_dfm_8) & mul_mul_mul_mul_nor_6_m1c
      & (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign MulIn_data_and_1_cse = core_wen & and_18_tmp;
  assign IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse = and_dcpl_38 | and_dcpl_39;
  assign else_MulOp_data_and_8_cse = core_wen & and_18_tmp & (~ mux_7_itm);
  assign or_27_cse = (cfg_precision!=2'b10);
  assign FpMul_8U_23U_oelse_1_and_4_cse = core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse
      & (~ mux_7_itm);
  assign else_MulOp_data_and_9_cse = core_wen & and_18_tmp & (~ mux_12_itm);
  assign FpMul_8U_23U_oelse_1_and_5_cse = core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse
      & (~ mux_12_itm);
  assign else_MulOp_data_and_10_cse = core_wen & and_18_tmp & (~ mux_17_itm);
  assign FpMul_8U_23U_oelse_1_and_6_cse = core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse
      & (~ mux_17_itm);
  assign else_MulOp_data_and_11_cse = core_wen & and_18_tmp & (~ mux_22_itm);
  assign FpMul_8U_23U_oelse_1_and_7_cse = core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse
      & (~ mux_22_itm);
  assign mul_mul_aelse_and_cse = core_wen & and_18_tmp & (~ io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign mux_26_nl = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_74_cse);
  assign MulIn_data_and_2_cse = core_wen & (~ and_dcpl_23) & (mux_26_nl);
  assign or_74_cse = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt;
  assign nor_319_nl = ~((~ main_stage_v_2) | mul_mul_land_1_lpi_1_dfm_5 | or_tmp_59);
  assign nor_320_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_6
      | mul_mul_land_1_lpi_1_dfm_st_5);
  assign mux_27_nl = MUX_s_1_2_2((nor_320_nl), (nor_319_nl), or_74_cse);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse = core_wen & (~ and_dcpl_23)
      & (mux_27_nl);
  assign nor_315_nl = ~((~ main_stage_v_2) | mul_mul_land_2_lpi_1_dfm_5 | or_tmp_75);
  assign nor_316_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_6
      | mul_mul_land_2_lpi_1_dfm_st_5);
  assign mux_29_nl = MUX_s_1_2_2((nor_316_nl), (nor_315_nl), or_74_cse);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse = core_wen & (~ and_dcpl_23)
      & (mux_29_nl);
  assign nor_311_nl = ~((~ main_stage_v_2) | mul_mul_land_3_lpi_1_dfm_5 | or_tmp_91);
  assign nor_312_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_6
      | mul_mul_land_3_lpi_1_dfm_st_5);
  assign mux_31_nl = MUX_s_1_2_2((nor_312_nl), (nor_311_nl), or_74_cse);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse = core_wen & (~ and_dcpl_23)
      & (mux_31_nl);
  assign nor_307_nl = ~((~ main_stage_v_2) | mul_mul_land_lpi_1_dfm_5 | or_tmp_107);
  assign nor_308_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_lpi_1_dfm_6
      | mul_mul_land_lpi_1_dfm_st_5);
  assign mux_33_nl = MUX_s_1_2_2((nor_308_nl), (nor_307_nl), or_74_cse);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse = core_wen & (~ and_dcpl_23)
      & (mux_33_nl);
  assign nor_20_cse = ~((cfg_precision!=2'b10));
  assign nor_301_cse = ~(FpMul_8U_23U_lor_6_lpi_1_dfm_6 | (~ (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1);
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse = and_dcpl_46 | and_dcpl_48
      | and_dcpl_50 | and_dcpl_51;
  assign FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse = and_dcpl_52
      | and_dcpl_47;
  assign nand_48_cse = ~(mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_2);
  assign IsNaN_8U_23U_1_aelse_and_cse = core_wen & (~ and_dcpl_23) & not_tmp_54;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse = MUX_s_1_2_2(mul_mul_1_FpMantRNE_48U_24U_else_and_tmp,
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st, and_dcpl_47);
  assign FpMantRNE_48U_24U_else_and_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_55;
  assign nor_277_cse = ~((~ (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1);
  assign nor_31_cse = ~(FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_282_cse = ~((~ mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2) | mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign IsNaN_8U_23U_aelse_and_17_cse = core_wen & (~ and_dcpl_23) & (~ mux_tmp_48);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_54;
  assign nor_264_cse = ~((~ (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | FpMul_8U_23U_lor_7_lpi_1_dfm_6);
  assign nor_348_cse = ~(FpMul_8U_23U_lor_7_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2);
  assign nor_267_cse = ~(nor_348_cse | mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse = and_dcpl_54 | and_dcpl_55
      | and_dcpl_57 | and_dcpl_58;
  assign nand_45_cse = ~(mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_2);
  assign IsNaN_8U_23U_1_aelse_and_1_cse = core_wen & (~ and_dcpl_23) & not_tmp_81;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse = MUX_s_1_2_2(mul_mul_2_FpMantRNE_48U_24U_else_and_tmp,
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st, and_dcpl_47);
  assign FpMantRNE_48U_24U_else_and_9_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_82;
  assign nor_241_cse = ~((~ (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1);
  assign nor_49_cse = ~(FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_245_cse = ~((~ mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2) | mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign IsNaN_8U_23U_aelse_and_19_cse = core_wen & (~ and_dcpl_23) & (~ mux_94_itm);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_81;
  assign nor_227_cse = ~((~ (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | FpMul_8U_23U_lor_8_lpi_1_dfm_6);
  assign nor_347_cse = ~(FpMul_8U_23U_lor_8_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2);
  assign nor_230_cse = ~(nor_347_cse | mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse = and_dcpl_60 | and_dcpl_61
      | and_dcpl_63 | and_dcpl_64;
  assign nand_42_cse = ~(mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_2);
  assign IsNaN_8U_23U_1_aelse_and_2_cse = core_wen & (~ and_dcpl_23) & not_tmp_106;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse = MUX_s_1_2_2(mul_mul_3_FpMantRNE_48U_24U_else_and_tmp,
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st, and_dcpl_47);
  assign FpMantRNE_48U_24U_else_and_11_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_107;
  assign nor_204_cse = ~((~ (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1);
  assign nor_68_cse = ~(FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_208_cse = ~((~ mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2) | mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign IsNaN_8U_23U_aelse_and_21_cse = core_wen & (~ and_dcpl_23) & (~ mux_125_itm);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_106;
  assign nor_190_cse = ~((~ (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | FpMul_8U_23U_lor_1_lpi_1_dfm_6);
  assign nor_346_cse = ~(FpMul_8U_23U_lor_1_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2);
  assign nor_193_cse = ~(nor_346_cse | mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2);
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse = and_dcpl_66 | and_dcpl_67
      | and_dcpl_69 | and_dcpl_70;
  assign or_430_cse = (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign IsNaN_8U_23U_1_aelse_and_3_cse = core_wen & (~ and_dcpl_23) & not_tmp_129;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse = MUX_s_1_2_2(mul_mul_4_FpMantRNE_48U_24U_else_and_tmp,
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st, and_dcpl_47);
  assign FpMantRNE_48U_24U_else_and_13_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_130;
  assign nor_170_cse = ~((~ (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1);
  assign nor_86_cse = ~(FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3));
  assign nor_174_cse = ~((~ mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2) | mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign IsNaN_8U_23U_aelse_and_23_cse = core_wen & (~ and_dcpl_23) & (~ mux_tmp_140);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse = core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
      & not_tmp_129;
  assign mul_mul_aelse_and_12_cse = core_wen & (~ and_dcpl_23) & (~ mux_tmp_46);
  assign MulIn_data_and_cse = core_wen & (~((~ and_20_tmp) | (fsm_output[0])));
  assign IsNaN_8U_23U_aelse_and_cse = core_wen & (~ (fsm_output[0]));
  assign IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse = and_dcpl_3 | and_dcpl_6;
  assign or_467_nl = mul_mul_land_1_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d;
  assign mux_160_nl = MUX_s_1_2_2(or_tmp_1, (or_467_nl), and_20_tmp);
  assign IsNaN_8U_23U_aelse_and_24_cse = IsNaN_8U_23U_aelse_and_cse & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse
      & (~ (mux_160_nl));
  assign or_480_nl = mul_mul_land_2_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d;
  assign mux_168_nl = MUX_s_1_2_2(or_tmp_15, (or_480_nl), and_20_tmp);
  assign IsNaN_8U_23U_aelse_and_25_cse = IsNaN_8U_23U_aelse_and_cse & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse
      & (~ (mux_168_nl));
  assign or_488_nl = mul_mul_land_3_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d;
  assign mux_173_nl = MUX_s_1_2_2(or_tmp_29, (or_488_nl), and_20_tmp);
  assign IsNaN_8U_23U_aelse_and_26_cse = IsNaN_8U_23U_aelse_and_cse & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse
      & (~ (mux_173_nl));
  assign or_496_nl = mul_mul_land_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d;
  assign mux_178_nl = MUX_s_1_2_2(or_tmp_46, (or_496_nl), and_20_tmp);
  assign IsNaN_8U_23U_aelse_and_27_cse = IsNaN_8U_23U_aelse_and_cse & IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse
      & (~ (mux_178_nl));
  assign mul_mul_aelse_and_19_cse = IsNaN_8U_23U_aelse_and_cse & and_20_tmp & (~
      cfg_mul_bypass_rsci_d);
  assign nor_143_cse = ~((~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt);
  assign FpMul_8U_23U_p_expo_and_cse = core_wen & (~ or_dcpl_22);
  assign else_MulOp_data_and_1_cse = core_wen & (~ or_dcpl_27);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_cse = core_wen & (~(or_dcpl_26
      | and_dcpl_37 | mul_mul_land_1_lpi_1_dfm_st_4));
  assign FpMul_8U_23U_p_expo_and_1_cse = core_wen & (~ or_dcpl_37);
  assign else_MulOp_data_and_3_cse = core_wen & (~ or_dcpl_40);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse = core_wen & (~(or_dcpl_26
      | and_dcpl_37 | mul_mul_land_2_lpi_1_dfm_st_4));
  assign FpMul_8U_23U_p_expo_and_2_cse = core_wen & (~ or_dcpl_50);
  assign else_MulOp_data_and_5_cse = core_wen & (~ or_dcpl_53);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse = core_wen & (~(or_dcpl_26
      | and_dcpl_37 | mul_mul_land_3_lpi_1_dfm_st_4));
  assign FpMul_8U_23U_p_expo_and_3_cse = core_wen & (~ or_dcpl_63);
  assign else_MulOp_data_and_7_cse = core_wen & (~ or_dcpl_66);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse = core_wen & (~(or_dcpl_26
      | and_dcpl_37 | mul_mul_land_lpi_1_dfm_st_4));
  assign and_136_m1c = and_18_tmp & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_4);
  assign and_135_rgt = and_18_tmp & IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  assign mul_mul_if_and_6_rgt = (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0) & and_136_m1c;
  assign mul_mul_if_and_7_rgt = IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 & and_136_m1c;
  assign and_138_m1c = and_18_tmp & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_4);
  assign and_137_rgt = and_18_tmp & IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  assign mul_mul_if_and_4_rgt = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0) & and_138_m1c;
  assign mul_mul_if_and_5_rgt = IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 & and_138_m1c;
  assign and_140_m1c = and_18_tmp & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_4);
  assign and_139_rgt = and_18_tmp & IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  assign mul_mul_if_and_2_rgt = (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0) & and_140_m1c;
  assign mul_mul_if_and_3_rgt = IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 & and_140_m1c;
  assign and_142_m1c = and_18_tmp & (~ IsNaN_8U_23U_land_lpi_1_dfm_4);
  assign and_141_rgt = and_18_tmp & IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign mul_mul_if_and_rgt = (~ IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0) & and_142_m1c;
  assign mul_mul_if_and_1_rgt = IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 & and_142_m1c;
  assign nor_118_cse = ~(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp | mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_land_1_lpi_1_dfm_4);
  assign and_146_rgt = (or_dcpl_75 | IsZero_8U_23U_land_1_lpi_1_dfm_4 | or_27_cse)
      & and_18_tmp;
  assign nor_117_cse = ~(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp | mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_land_2_lpi_1_dfm_4);
  assign and_150_rgt = (or_dcpl_81 | IsZero_8U_23U_land_2_lpi_1_dfm_4 | or_27_cse)
      & and_18_tmp;
  assign nor_116_cse = ~(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp | mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_land_3_lpi_1_dfm_4);
  assign and_154_rgt = (or_dcpl_87 | IsZero_8U_23U_land_3_lpi_1_dfm_4 | or_27_cse)
      & and_18_tmp;
  assign nor_115_cse = ~(IsZero_8U_23U_land_lpi_1_dfm_4 | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp
      | mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1);
  assign and_158_rgt = (or_dcpl_93 | mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 |
      or_27_cse) & and_18_tmp;
  assign or_468_cse = (~ and_18_tmp) | (cfg_precision!=2'b10);
  assign or_469_cse = (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs)
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st;
  assign or_482_cse = (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs)
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st;
  assign or_490_cse = (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs)
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st;
  assign IsNaN_8U_23U_aelse_and_4_cse = core_wen & (~((cfg_mul_prelu_rsci_d & (~
      (chn_mul_in_rsci_d_mxwt[31]))) | cfg_mul_bypass_rsci_d | or_dcpl_110 | (fsm_output[0])));
  assign IsNaN_8U_23U_aelse_and_5_cse = core_wen & (~((cfg_mul_prelu_rsci_d & (~
      (chn_mul_in_rsci_d_mxwt[63]))) | cfg_mul_bypass_rsci_d | or_dcpl_110 | (fsm_output[0])));
  assign IsNaN_8U_23U_aelse_and_6_cse = core_wen & (~((cfg_mul_prelu_rsci_d & (~
      (chn_mul_in_rsci_d_mxwt[95]))) | cfg_mul_bypass_rsci_d | or_dcpl_110 | (fsm_output[0])));
  assign IsNaN_8U_23U_aelse_and_7_cse = core_wen & (~((cfg_mul_prelu_rsci_d & (~
      (chn_mul_in_rsci_d_mxwt[127]))) | cfg_mul_bypass_rsci_d | or_dcpl_110 | (fsm_output[0])));
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp = ~((else_MulOp_data_0_lpi_1_dfm_mx0_30_0!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp = ~((else_MulOp_data_1_lpi_1_dfm_mx0_30_0!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp = ~((else_MulOp_data_2_lpi_1_dfm_mx0_30_0!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp = ~((else_MulOp_data_3_lpi_1_dfm_mx0_30_0!=31'b0000000000000000000000000000000));
  assign nl_FpMul_8U_23U_else_2_else_acc_nl = (else_MulOp_data_0_lpi_1_dfm_2_30_0_1[30:23])
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_nl = nl_FpMul_8U_23U_else_2_else_acc_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_nl)
      + (MulIn_data_sva_132[30:23]);
  assign FpMul_8U_23U_p_expo_1_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0 = ~(mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      & (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_mul_1_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_1_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_1_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_1_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_1_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0 = (mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | (~ (FpMul_8U_23U_p_mant_p1_1_sva_mx1[47]))) & mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[63:31]==33'b111111111111111111111111111111111));
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[63:31]!=33'b000000000000000000000000000000000));
  assign nl_FpMul_8U_23U_else_2_else_acc_2_nl = (else_MulOp_data_1_lpi_1_dfm_2_30_0_1[30:23])
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_2_nl = nl_FpMul_8U_23U_else_2_else_acc_2_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_2_nl)
      + (MulIn_data_sva_132[62:55]);
  assign FpMul_8U_23U_p_expo_2_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0 = ~(mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      & (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_mul_2_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_2_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_2_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_2_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_2_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0 = (mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | (~ (FpMul_8U_23U_p_mant_p1_2_sva_mx1[47]))) & mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[63:31]==33'b111111111111111111111111111111111));
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[63:31]!=33'b000000000000000000000000000000000));
  assign nl_FpMul_8U_23U_else_2_else_acc_3_nl = (else_MulOp_data_2_lpi_1_dfm_2_30_0_1[30:23])
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_3_nl = nl_FpMul_8U_23U_else_2_else_acc_3_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_3_nl)
      + (MulIn_data_sva_132[94:87]);
  assign FpMul_8U_23U_p_expo_3_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0 = ~(mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      & (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_mul_3_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_3_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_3_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_3_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_3_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0 = (mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | (~ (FpMul_8U_23U_p_mant_p1_3_sva_mx1[47]))) & mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[63:31]==33'b111111111111111111111111111111111));
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[63:31]!=33'b000000000000000000000000000000000));
  assign nl_FpMul_8U_23U_else_2_else_acc_4_nl = (else_MulOp_data_3_lpi_1_dfm_2_30_0_1[30:23])
      + 8'b10000001;
  assign FpMul_8U_23U_else_2_else_acc_4_nl = nl_FpMul_8U_23U_else_2_else_acc_4_nl[7:0];
  assign nl_FpMul_8U_23U_p_expo_sva_1_mx0w0 = (FpMul_8U_23U_else_2_else_acc_4_nl)
      + (MulIn_data_sva_132[126:119]);
  assign FpMul_8U_23U_p_expo_sva_1_mx0w0 = nl_FpMul_8U_23U_p_expo_sva_1_mx0w0[7:0];
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0 = ~(mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      & (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]));
  assign mul_mul_4_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_sva_mx0w0
      & (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23]==23'b11111111111111111111111);
  assign FpMantRNE_48U_24U_else_carry_sva_mx0w0 = (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[22])
      & (((FpMul_8U_23U_p_mant_p1_sva_mx1[0]) & (FpMul_8U_23U_p_mant_p1_sva_mx1[47]))
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[0]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[2]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[4]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[6]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[8]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[9])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[10]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[11])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[12]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[13])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[14]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[15])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[16]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[17])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[18]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[19])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[20]) | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[21])
      | (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[23]));
  assign FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0 = (mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1
      | (~ (FpMul_8U_23U_p_mant_p1_sva_mx1[47]))) & mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[63:31]==33'b111111111111111111111111111111111));
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[63:31]!=33'b000000000000000000000000000000000));
  assign IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[62:32]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[94:64]!=31'b0000000000000000000000000000000));
  assign IsZero_8U_23U_land_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[126:96]!=31'b0000000000000000000000000000000));
  assign mul_mul_land_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[127]) | (~ cfg_mul_prelu_rsci_d));
  assign mul_mul_land_3_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[95]) | (~ cfg_mul_prelu_rsci_d));
  assign mul_mul_land_2_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[63]) | (~ cfg_mul_prelu_rsci_d));
  assign mul_mul_land_1_lpi_1_dfm_mx1w0 = ~((chn_mul_in_rsci_d_mxwt[31]) | (~ cfg_mul_prelu_rsci_d));
  assign FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 = mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp | IsZero_8U_23U_land_1_lpi_1_dfm_4;
  assign IsNaN_8U_23U_1_nor_tmp = ~((else_MulOp_data_0_lpi_1_dfm_mx0_30_0[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_1_nor_tmp | (else_MulOp_data_0_lpi_1_dfm_mx0_30_0[30:23]!=8'b11111111));
  assign FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0 = mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp | IsZero_8U_23U_land_2_lpi_1_dfm_4;
  assign IsNaN_8U_23U_1_nor_1_tmp = ~((else_MulOp_data_1_lpi_1_dfm_mx0_30_0[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_1_nor_1_tmp | (else_MulOp_data_1_lpi_1_dfm_mx0_30_0[30:23]!=8'b11111111));
  assign FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 = mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp | IsZero_8U_23U_land_3_lpi_1_dfm_4;
  assign IsNaN_8U_23U_1_nor_2_tmp = ~((else_MulOp_data_2_lpi_1_dfm_mx0_30_0[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_1_nor_2_tmp | (else_MulOp_data_2_lpi_1_dfm_mx0_30_0[30:23]!=8'b11111111));
  assign FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0 = mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp | IsZero_8U_23U_land_lpi_1_dfm_4;
  assign IsNaN_8U_23U_1_nor_3_tmp = ~((else_MulOp_data_3_lpi_1_dfm_mx0_30_0[22:0]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_1_nor_3_tmp | (else_MulOp_data_3_lpi_1_dfm_mx0_30_0[30:23]!=8'b11111111));
  assign FpMul_8U_23U_p_mant_p1_and_7_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_6_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_1_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_1_sva,
      mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_7_nl);
  assign mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_1_lpi_1_dfm_6)
      , (MulIn_data_sva_132[22:0])}) * ({(~ IsZero_8U_23U_1_land_1_lpi_1_dfm_6) ,
      (else_MulOp_data_0_lpi_1_dfm_2_30_0_1[22:0])}));
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_1[30:23])
      + conv_u2u_8_9(else_MulOp_data_0_lpi_1_dfm_mx0_30_0[30:23]);
  assign mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl));
  assign mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = conv_s2u_64_64($signed((MulIn_data_sva_1[31:0]))
      * $signed(else_MulOp_data_0_lpi_1_dfm_mx1));
  assign FpMul_8U_23U_p_mant_p1_and_6_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_7_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_2_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_2_sva,
      mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_6_nl);
  assign mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_2_lpi_1_dfm_6)
      , (MulIn_data_sva_132[54:32])}) * ({(~ IsZero_8U_23U_1_land_2_lpi_1_dfm_6)
      , (else_MulOp_data_1_lpi_1_dfm_2_30_0_1[22:0])}));
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_1[62:55])
      + conv_u2u_8_9(else_MulOp_data_1_lpi_1_dfm_mx0_30_0[30:23]);
  assign mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl));
  assign mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = conv_s2u_64_64($signed((MulIn_data_sva_1[63:32]))
      * $signed(else_MulOp_data_1_lpi_1_dfm_mx1));
  assign FpMul_8U_23U_p_mant_p1_and_5_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_8_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_3_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_3_sva,
      mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_5_nl);
  assign mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_3_lpi_1_dfm_6)
      , (MulIn_data_sva_132[86:64])}) * ({(~ IsZero_8U_23U_1_land_3_lpi_1_dfm_6)
      , (else_MulOp_data_2_lpi_1_dfm_2_30_0_1[22:0])}));
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_1[94:87])
      + conv_u2u_8_9(else_MulOp_data_2_lpi_1_dfm_mx0_30_0[30:23]);
  assign mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl));
  assign mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = conv_s2u_64_64($signed((MulIn_data_sva_1[95:64]))
      * $signed(else_MulOp_data_2_lpi_1_dfm_mx1));
  assign FpMul_8U_23U_p_mant_p1_and_4_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & (~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_3);
  assign FpMul_8U_23U_p_mant_p1_sva_mx1 = MUX_v_48_2_2(FpMul_8U_23U_p_mant_p1_sva,
      mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp, FpMul_8U_23U_p_mant_p1_and_4_nl);
  assign mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp = conv_u2u_48_48(({(~ IsZero_8U_23U_land_lpi_1_dfm_6)
      , (MulIn_data_sva_132[118:96])}) * ({(~ IsZero_8U_23U_1_land_lpi_1_dfm_6) ,
      (else_MulOp_data_3_lpi_1_dfm_2_30_0_1[22:0])}));
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl = conv_u2u_8_9(MulIn_data_sva_1[126:119])
      + conv_u2u_8_9(else_MulOp_data_3_lpi_1_dfm_mx0_30_0[30:23]);
  assign mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl = nl_mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl[8:0];
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl = conv_u2u_8_9(readslicef_9_8_1((mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl)))
      + 9'b101000001;
  assign mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl = nl_mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8:0];
  assign mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1 = readslicef_9_1_8((mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl));
  assign mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = conv_s2u_64_64($signed((MulIn_data_sva_1[127:96]))
      * $signed(else_MulOp_data_3_lpi_1_dfm_mx1));
  assign IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[62:55]!=8'b11111111));
  assign IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[94:87]!=8'b11111111));
  assign IsNaN_8U_23U_land_lpi_1_dfm_mx0w0 = ~((~((chn_mul_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000)))
      | (chn_mul_in_rsci_d_mxwt[126:119]!=8'b11111111));
  assign nl_mul_mul_1_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_1_sva_2);
  assign mul_mul_1_FpMantRNE_48U_24U_else_acc_nl = nl_mul_mul_1_FpMantRNE_48U_24U_else_acc_nl[22:0];
  assign or_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp | (~ mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2);
  assign mux_237_nl = MUX_v_23_2_2((signext_23_1(~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp)),
      (mul_mul_1_FpMantRNE_48U_24U_else_acc_nl), or_nl);
  assign FpMul_8U_23U_nor_nl = ~(MUX_v_23_2_2((mux_237_nl), 23'b11111111111111111111111,
      FpMul_8U_23U_is_inf_1_lpi_1_dfm_2));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_4_nl = ~(MUX_v_23_2_2((FpMul_8U_23U_nor_nl),
      23'b11111111111111111111111, FpMul_8U_23U_lor_9_lpi_1_dfm));
  assign FpMul_8U_23U_FpMul_8U_23U_nor_nl = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 |
      IsNaN_8U_23U_land_1_lpi_1_dfm_8);
  assign FpMul_8U_23U_and_1_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_8);
  assign FpMul_8U_23U_o_mant_1_lpi_1_dfm_3 = MUX1HOT_v_23_3_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_4_nl),
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2, (MulIn_data_sva_133[22:0]),
      {(FpMul_8U_23U_FpMul_8U_23U_nor_nl) , (FpMul_8U_23U_and_1_nl) , IsNaN_8U_23U_land_1_lpi_1_dfm_8});
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva = ~(IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1
      | mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1
      & mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign mul_mul_else_unequal_tmp_1 = ~((cfg_precision==2'b10));
  assign nl_mul_mul_2_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_2_sva_2);
  assign mul_mul_2_FpMantRNE_48U_24U_else_acc_nl = nl_mul_mul_2_FpMantRNE_48U_24U_else_acc_nl[22:0];
  assign or_840_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1 | (~ mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2);
  assign mux_238_nl = MUX_v_23_2_2((signext_23_1(~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1)),
      (mul_mul_2_FpMantRNE_48U_24U_else_acc_nl), or_840_nl);
  assign FpMul_8U_23U_nor_4_nl = ~(MUX_v_23_2_2((mux_238_nl), 23'b11111111111111111111111,
      nor_348_cse));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_5_nl = ~(MUX_v_23_2_2((FpMul_8U_23U_nor_4_nl),
      23'b11111111111111111111111, FpMul_8U_23U_lor_10_lpi_1_dfm));
  assign FpMul_8U_23U_FpMul_8U_23U_nor_1_nl = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      | IsNaN_8U_23U_land_2_lpi_1_dfm_8);
  assign FpMul_8U_23U_and_3_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_8);
  assign FpMul_8U_23U_o_mant_2_lpi_1_dfm_3 = MUX1HOT_v_23_3_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_5_nl),
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2, (MulIn_data_sva_133[54:32]),
      {(FpMul_8U_23U_FpMul_8U_23U_nor_1_nl) , (FpMul_8U_23U_and_3_nl) , IsNaN_8U_23U_land_2_lpi_1_dfm_8});
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva = ~(IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1
      | mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1
      & mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign nl_mul_mul_3_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_3_sva_2);
  assign mul_mul_3_FpMantRNE_48U_24U_else_acc_nl = nl_mul_mul_3_FpMantRNE_48U_24U_else_acc_nl[22:0];
  assign or_841_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2 | (~ mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2);
  assign mux_239_nl = MUX_v_23_2_2((signext_23_1(~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2)),
      (mul_mul_3_FpMantRNE_48U_24U_else_acc_nl), or_841_nl);
  assign FpMul_8U_23U_nor_5_nl = ~(MUX_v_23_2_2((mux_239_nl), 23'b11111111111111111111111,
      nor_347_cse));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_6_nl = ~(MUX_v_23_2_2((FpMul_8U_23U_nor_5_nl),
      23'b11111111111111111111111, FpMul_8U_23U_lor_11_lpi_1_dfm));
  assign FpMul_8U_23U_FpMul_8U_23U_nor_2_nl = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      | IsNaN_8U_23U_land_3_lpi_1_dfm_8);
  assign FpMul_8U_23U_and_5_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_8);
  assign FpMul_8U_23U_o_mant_3_lpi_1_dfm_3 = MUX1HOT_v_23_3_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_6_nl),
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2, (MulIn_data_sva_133[86:64]),
      {(FpMul_8U_23U_FpMul_8U_23U_nor_2_nl) , (FpMul_8U_23U_and_5_nl) , IsNaN_8U_23U_land_3_lpi_1_dfm_8});
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva = ~(IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1
      | mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1
      & mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign nl_mul_mul_4_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2
      + conv_u2u_1_23(FpMantRNE_48U_24U_else_carry_sva_2);
  assign mul_mul_4_FpMantRNE_48U_24U_else_acc_nl = nl_mul_mul_4_FpMantRNE_48U_24U_else_acc_nl[22:0];
  assign or_842_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3 | (~ mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2);
  assign mux_240_nl = MUX_v_23_2_2((signext_23_1(~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3)),
      (mul_mul_4_FpMantRNE_48U_24U_else_acc_nl), or_842_nl);
  assign FpMul_8U_23U_nor_6_nl = ~(MUX_v_23_2_2((mux_240_nl), 23'b11111111111111111111111,
      nor_346_cse));
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_7_nl = ~(MUX_v_23_2_2((FpMul_8U_23U_nor_6_nl),
      23'b11111111111111111111111, FpMul_8U_23U_lor_2_lpi_1_dfm));
  assign FpMul_8U_23U_FpMul_8U_23U_nor_3_nl = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_7 |
      IsNaN_8U_23U_land_lpi_1_dfm_8);
  assign FpMul_8U_23U_and_7_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & (~ IsNaN_8U_23U_land_lpi_1_dfm_8);
  assign FpMul_8U_23U_o_mant_lpi_1_dfm_3 = MUX1HOT_v_23_3_2((FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_7_nl),
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2, (MulIn_data_sva_133[118:96]),
      {(FpMul_8U_23U_FpMul_8U_23U_nor_3_nl) , (FpMul_8U_23U_and_7_nl) , IsNaN_8U_23U_land_lpi_1_dfm_8});
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva = ~(IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1
      | mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2);
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1
      & mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign mul_mul_mul_mul_nor_6_m1c = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_lpi_1_dfm_6);
  assign mul_mul_mul_mul_nor_4_m1c = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_3_lpi_1_dfm_6);
  assign mul_mul_mul_mul_nor_2_m1c = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_2_lpi_1_dfm_6);
  assign mul_mul_mul_mul_nor_m1c = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_1_lpi_1_dfm_6);
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_1_sva_5
      + 8'b1;
  assign mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      FpMul_8U_23U_p_expo_1_sva_5, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 = FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1[7:0];
  assign FpMul_8U_23U_FpMul_8U_23U_nor_4_nl = ~(mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2
      | FpMul_8U_23U_is_inf_1_lpi_1_dfm_2);
  assign FpMul_8U_23U_or_4_nl = ((~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp)
      & mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2) | FpMul_8U_23U_is_inf_1_lpi_1_dfm_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp
      & mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2 & (~ FpMul_8U_23U_is_inf_1_lpi_1_dfm_2);
  assign FpMul_8U_23U_o_expo_1_lpi_1_dfm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1, {(FpMul_8U_23U_FpMul_8U_23U_nor_4_nl)
      , (FpMul_8U_23U_or_4_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl)});
  assign FpMul_8U_23U_lor_9_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_1_lpi_1_dfm!=8'b00000000)))
      | FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  assign FpMul_8U_23U_is_inf_1_lpi_1_dfm_2 = ~(FpMul_8U_23U_FpMul_8U_23U_and_itm_2
      | FpMul_8U_23U_lor_6_lpi_1_dfm_7);
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_2_sva_5
      + 8'b1;
  assign mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      FpMul_8U_23U_p_expo_2_sva_5, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 = FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1[7:0];
  assign FpMul_8U_23U_or_5_nl = ((~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1)
      & mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2) | nor_348_cse;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1
      & mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2 & (~ nor_348_cse);
  assign FpMul_8U_23U_o_expo_2_lpi_1_dfm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1, {nor_267_cse ,
      (FpMul_8U_23U_or_5_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl)});
  assign FpMul_8U_23U_lor_10_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_2_lpi_1_dfm!=8'b00000000)))
      | FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_3_sva_5
      + 8'b1;
  assign mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      FpMul_8U_23U_p_expo_3_sva_5, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 = FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1[7:0];
  assign FpMul_8U_23U_or_6_nl = ((~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2)
      & mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2) | nor_347_cse;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2
      & mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2 & (~ nor_347_cse);
  assign FpMul_8U_23U_o_expo_3_lpi_1_dfm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1, {nor_230_cse ,
      (FpMul_8U_23U_or_6_nl) , (FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl)});
  assign FpMul_8U_23U_lor_11_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_3_lpi_1_dfm!=8'b00000000)))
      | FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_sva_5
      + 8'b1;
  assign mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl = nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0];
  assign FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl),
      FpMul_8U_23U_p_expo_sva_5, FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2);
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3 = ~((FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1==8'b11111111));
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0
      + 8'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1[7:0];
  assign FpMul_8U_23U_or_7_nl = ((~ FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3)
      & mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2) | nor_346_cse;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3
      & mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2 & (~ nor_346_cse);
  assign FpMul_8U_23U_o_expo_lpi_1_dfm = MUX1HOT_v_8_3_2(FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0,
      8'b11111110, FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1, {nor_193_cse , (FpMul_8U_23U_or_7_nl)
      , (FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl)});
  assign FpMul_8U_23U_lor_2_lpi_1_dfm = (~((FpMul_8U_23U_o_expo_lpi_1_dfm!=8'b00000000)))
      | FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  assign nl_FpMul_8U_23U_oelse_1_acc_nl = conv_u2s_8_9(else_MulOp_data_0_lpi_1_dfm_mx0_30_0[30:23])
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_nl = nl_FpMul_8U_23U_oelse_1_acc_nl[8:0];
  assign nl_mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_nl)
      + conv_u2s_8_10(MulIn_data_sva_1[30:23]);
  assign mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl));
  assign else_MulOp_data_0_lpi_1_dfm_mx0_30_0 = MUX_v_31_2_2((cfg_mul_op_1_sva_1[30:0]),
      (chn_mul_op_rsci_d_mxwt[30:0]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_0_lpi_1_dfm_mx1 = MUX_v_32_2_2(cfg_mul_op_1_sva_1, (chn_mul_op_rsci_d_mxwt[31:0]),
      cfg_mul_src_1_sva_1);
  assign nl_FpMul_8U_23U_oelse_1_acc_1_nl = conv_u2s_8_9(else_MulOp_data_1_lpi_1_dfm_mx0_30_0[30:23])
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_1_nl = nl_FpMul_8U_23U_oelse_1_acc_1_nl[8:0];
  assign nl_mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_1_nl)
      + conv_u2s_8_10(MulIn_data_sva_1[62:55]);
  assign mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl));
  assign else_MulOp_data_1_lpi_1_dfm_mx0_30_0 = MUX_v_31_2_2((cfg_mul_op_1_sva_1[30:0]),
      (chn_mul_op_rsci_d_mxwt[62:32]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_1_lpi_1_dfm_mx1 = MUX_v_32_2_2(cfg_mul_op_1_sva_1, (chn_mul_op_rsci_d_mxwt[63:32]),
      cfg_mul_src_1_sva_1);
  assign nl_FpMul_8U_23U_oelse_1_acc_2_nl = conv_u2s_8_9(else_MulOp_data_2_lpi_1_dfm_mx0_30_0[30:23])
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_2_nl = nl_FpMul_8U_23U_oelse_1_acc_2_nl[8:0];
  assign nl_mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_2_nl)
      + conv_u2s_8_10(MulIn_data_sva_1[94:87]);
  assign mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl));
  assign else_MulOp_data_2_lpi_1_dfm_mx0_30_0 = MUX_v_31_2_2((cfg_mul_op_1_sva_1[30:0]),
      (chn_mul_op_rsci_d_mxwt[94:64]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_2_lpi_1_dfm_mx1 = MUX_v_32_2_2(cfg_mul_op_1_sva_1, (chn_mul_op_rsci_d_mxwt[95:64]),
      cfg_mul_src_1_sva_1);
  assign nl_FpMul_8U_23U_oelse_1_acc_3_nl = conv_u2s_8_9(else_MulOp_data_3_lpi_1_dfm_mx0_30_0[30:23])
      + 9'b110000001;
  assign FpMul_8U_23U_oelse_1_acc_3_nl = nl_FpMul_8U_23U_oelse_1_acc_3_nl[8:0];
  assign nl_mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl = conv_s2s_9_10(FpMul_8U_23U_oelse_1_acc_3_nl)
      + conv_u2s_8_10(MulIn_data_sva_1[126:119]);
  assign mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl = nl_mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9:0];
  assign mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 = readslicef_10_1_9((mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl));
  assign else_MulOp_data_3_lpi_1_dfm_mx0_30_0 = MUX_v_31_2_2((cfg_mul_op_1_sva_1[30:0]),
      (chn_mul_op_rsci_d_mxwt[126:96]), cfg_mul_src_1_sva_1);
  assign else_MulOp_data_3_lpi_1_dfm_mx1 = MUX_v_32_2_2(cfg_mul_op_1_sva_1, (chn_mul_op_rsci_d_mxwt[127:96]),
      cfg_mul_src_1_sva_1);
  assign and_20_tmp = chn_mul_in_rsci_bawt & or_11_cse & or_12_cse & or_13_cse &
      or_14_cse & or_15_cse & or_16_cse & or_74_cse;
  assign or_11_cse = chn_mul_op_rsci_bawt | (~(cfg_mul_src_1_sva_st_1 & (~ io_read_cfg_mul_bypass_rsc_svs_st_1)
      & main_stage_v_1));
  assign or_12_cse = cfg_truncate_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_13_cse = cfg_mul_op_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_14_cse = cfg_mul_src_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_15_cse = cfg_mul_prelu_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign or_16_cse = cfg_mul_bypass_rsc_triosy_obj_bawt | (~ main_stage_v_1);
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1022])
      & ((IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[0]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[2]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[3])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[4]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[5])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[6]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[7])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[8]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[9])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[10]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[11])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[12]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[13])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[14]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[15])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[16]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[17])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[18]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[19])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[20]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[21])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[22]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[23])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[24]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[25])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[26]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[27])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[28]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[29])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[30]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[31])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[32]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[33])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[34]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[35])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[36]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[37])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[38]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[39])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[40]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[41])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[42]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[43])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[44]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[45])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[46]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[47])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[48]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[49])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[50]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[51])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[52]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[53])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[54]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[55])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[56]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[57])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[58]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[59])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[60]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[61])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[62]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[63])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[64]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[65])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[66]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[67])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[68]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[69])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[70]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[71])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[72]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[73])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[74]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[75])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[76]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[77])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[78]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[79])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[80]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[81])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[82]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[83])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[84]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[85])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[86]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[87])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[88]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[89])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[90]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[91])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[92]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[93])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[94]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[95])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[96]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[97])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[98]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[99])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[100]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[101])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[102]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[103])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[104]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[105])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[106]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[107])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[108]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[109])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[110]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[111])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[112]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[113])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[114]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[115])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[116]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[117])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[118]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[119])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[120]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[121])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[122]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[123])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[124]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[125])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[126]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[127])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[128]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[129])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[130]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[131])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[132]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[133])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[134]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[135])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[136]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[137])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[138]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[139])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[140]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[141])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[142]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[143])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[144]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[145])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[146]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[147])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[148]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[149])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[150]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[151])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[152]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[153])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[154]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[155])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[156]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[157])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[158]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[159])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[160]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[161])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[162]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[163])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[164]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[165])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[166]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[167])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[168]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[169])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[170]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[171])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[172]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[173])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[174]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[175])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[176]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[177])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[178]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[179])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[180]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[181])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[182]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[183])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[184]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[185])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[186]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[187])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[188]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[189])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[190]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[191])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[192]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[193])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[194]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[195])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[196]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[197])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[198]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[199])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[200]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[201])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[202]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[203])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[204]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[205])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[206]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[207])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[208]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[209])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[210]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[211])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[212]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[213])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[214]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[215])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[216]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[217])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[218]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[219])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[220]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[221])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[222]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[223])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[224]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[225])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[226]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[227])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[228]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[229])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[230]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[231])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[232]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[233])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[234]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[235])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[236]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[237])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[238]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[239])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[240]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[241])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[242]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[243])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[244]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[245])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[246]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[247])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[248]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[249])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[250]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[251])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[252]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[253])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[254]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[255])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[256]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[257])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[258]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[259])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[260]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[261])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[262]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[263])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[264]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[265])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[266]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[267])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[268]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[269])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[270]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[271])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[272]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[273])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[274]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[275])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[276]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[277])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[278]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[279])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[280]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[281])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[282]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[283])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[284]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[285])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[286]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[287])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[288]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[289])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[290]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[291])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[292]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[293])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[294]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[295])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[296]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[297])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[298]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[299])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[300]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[301])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[302]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[303])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[304]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[305])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[306]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[307])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[308]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[309])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[310]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[311])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[312]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[313])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[314]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[315])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[316]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[317])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[318]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[319])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[320]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[321])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[322]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[323])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[324]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[325])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[326]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[327])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[328]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[329])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[330]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[331])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[332]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[333])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[334]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[335])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[336]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[337])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[338]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[339])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[340]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[341])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[342]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[343])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[344]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[345])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[346]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[347])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[348]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[349])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[350]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[351])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[352]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[353])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[354]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[355])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[356]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[357])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[358]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[359])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[360]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[361])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[362]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[363])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[364]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[365])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[366]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[367])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[368]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[369])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[370]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[371])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[372]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[373])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[374]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[375])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[376]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[377])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[378]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[379])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[380]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[381])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[382]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[383])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[384]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[385])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[386]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[387])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[388]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[389])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[390]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[391])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[392]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[393])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[394]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[395])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[396]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[397])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[398]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[399])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[400]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[401])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[402]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[403])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[404]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[405])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[406]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[407])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[408]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[409])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[410]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[411])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[412]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[413])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[414]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[415])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[416]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[417])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[418]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[419])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[420]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[421])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[422]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[423])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[424]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[425])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[426]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[427])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[428]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[429])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[430]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[431])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[432]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[433])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[434]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[435])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[436]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[437])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[438]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[439])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[440]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[441])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[442]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[443])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[444]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[445])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[446]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[447])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[448]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[449])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[450]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[451])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[452]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[453])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[454]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[455])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[456]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[457])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[458]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[459])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[460]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[461])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[462]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[463])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[464]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[465])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[466]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[467])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[468]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[469])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[470]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[471])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[472]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[473])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[474]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[475])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[476]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[477])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[478]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[479])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[480]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[481])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[482]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[483])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[484]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[485])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[486]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[487])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[488]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[489])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[490]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[491])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[492]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[493])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[494]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[495])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[496]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[497])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[498]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[499])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[500]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[501])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[502]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[503])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[504]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[505])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[506]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[507])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[508]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[509])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[510]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[511])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[512]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[513])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[514]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[515])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[516]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[517])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[518]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[519])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[520]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[521])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[522]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[523])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[524]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[525])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[526]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[527])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[528]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[529])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[530]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[531])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[532]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[533])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[534]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[535])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[536]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[537])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[538]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[539])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[540]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[541])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[542]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[543])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[544]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[545])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[546]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[547])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[548]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[549])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[550]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[551])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[552]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[553])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[554]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[555])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[556]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[557])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[558]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[559])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[560]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[561])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[562]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[563])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[564]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[565])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[566]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[567])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[568]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[569])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[570]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[571])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[572]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[573])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[574]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[575])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[576]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[577])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[578]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[579])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[580]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[581])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[582]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[583])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[584]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[585])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[586]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[587])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[588]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[589])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[590]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[591])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[592]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[593])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[594]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[595])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[596]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[597])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[598]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[599])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[600]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[601])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[602]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[603])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[604]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[605])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[606]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[607])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[608]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[609])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[610]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[611])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[612]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[613])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[614]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[615])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[616]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[617])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[618]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[619])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[620]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[621])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[622]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[623])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[624]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[625])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[626]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[627])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[628]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[629])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[630]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[631])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[632]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[633])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[634]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[635])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[636]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[637])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[638]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[639])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[640]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[641])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[642]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[643])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[644]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[645])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[646]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[647])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[648]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[649])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[650]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[651])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[652]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[653])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[654]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[655])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[656]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[657])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[658]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[659])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[660]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[661])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[662]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[663])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[664]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[665])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[666]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[667])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[668]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[669])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[670]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[671])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[672]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[673])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[674]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[675])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[676]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[677])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[678]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[679])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[680]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[681])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[682]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[683])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[684]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[685])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[686]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[687])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[688]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[689])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[690]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[691])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[692]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[693])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[694]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[695])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[696]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[697])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[698]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[699])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[700]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[701])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[702]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[703])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[704]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[705])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[706]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[707])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[708]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[709])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[710]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[711])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[712]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[713])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[714]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[715])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[716]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[717])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[718]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[719])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[720]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[721])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[722]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[723])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[724]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[725])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[726]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[727])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[728]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[729])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[730]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[731])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[732]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[733])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[734]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[735])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[736]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[737])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[738]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[739])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[740]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[741])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[742]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[743])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[744]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[745])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[746]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[747])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[748]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[749])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[750]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[751])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[752]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[753])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[754]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[755])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[756]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[757])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[758]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[759])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[760]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[761])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[762]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[763])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[764]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[765])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[766]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[767])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[768]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[769])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[770]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[771])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[772]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[773])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[774]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[775])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[776]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[777])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[778]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[779])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[780]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[781])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[782]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[783])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[784]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[785])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[786]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[787])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[788]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[789])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[790]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[791])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[792]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[793])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[794]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[795])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[796]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[797])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[798]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[799])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[800]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[801])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[802]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[803])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[804]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[805])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[806]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[807])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[808]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[809])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[810]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[811])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[812]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[813])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[814]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[815])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[816]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[817])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[818]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[819])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[820]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[821])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[822]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[823])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[824]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[825])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[826]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[827])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[828]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[829])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[830]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[831])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[832]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[833])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[834]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[835])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[836]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[837])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[838]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[839])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[840]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[841])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[842]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[843])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[844]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[845])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[846]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[847])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[848]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[849])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[850]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[851])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[852]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[853])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[854]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[855])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[856]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[857])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[858]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[859])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[860]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[861])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[862]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[863])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[864]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[865])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[866]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[867])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[868]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[869])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[870]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[871])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[872]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[873])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[874]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[875])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[876]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[877])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[878]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[879])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[880]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[881])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[882]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[883])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[884]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[885])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[886]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[887])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[888]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[889])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[890]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[891])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[892]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[893])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[894]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[895])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[896]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[897])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[898]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[899])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[900]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[901])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[902]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[903])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[904]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[905])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[906]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[907])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[908]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[909])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[910]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[911])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[912]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[913])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[914]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[915])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[916]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[917])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[918]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[919])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[920]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[921])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[922]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[923])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[924]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[925])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[926]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[927])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[928]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[929])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[930]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[931])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[932]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[933])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[934]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[935])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[936]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[937])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[938]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[939])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[940]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[941])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[942]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[943])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[944]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[945])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[946]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[947])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[948]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[949])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[950]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[951])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[952]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[953])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[954]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[955])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[956]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[957])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[958]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[959])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[960]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[961])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[962]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[963])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[964]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[965])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[966]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[967])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[968]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[969])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[970]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[971])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[972]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[973])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[974]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[975])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[976]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[977])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[978]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[979])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[980]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[981])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[982]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[983])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[984]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[985])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[986]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[987])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[988]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[989])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[990]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[991])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[992]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[993])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[994]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[995])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[996]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[997])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[998]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[999])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1000]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1001])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1002]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1003])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1004]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1005])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1006]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1007])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1008]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1009])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1010]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1011])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1012]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1013])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1014]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1015])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1016]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1017])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1018]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1019])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1020]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1021])
      | (~ (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1086])));
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva = conv_s2s_64_65(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1086:1023])
      + conv_u2s_1_65(mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_and_nl);
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva = nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[64:0];
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1022])
      & ((IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[0]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[2]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[3])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[4]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[5])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[6]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[7])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[8]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[9])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[10]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[11])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[12]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[13])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[14]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[15])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[16]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[17])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[18]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[19])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[20]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[21])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[22]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[23])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[24]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[25])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[26]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[27])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[28]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[29])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[30]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[31])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[32]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[33])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[34]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[35])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[36]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[37])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[38]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[39])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[40]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[41])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[42]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[43])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[44]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[45])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[46]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[47])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[48]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[49])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[50]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[51])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[52]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[53])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[54]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[55])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[56]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[57])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[58]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[59])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[60]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[61])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[62]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[63])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[64]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[65])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[66]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[67])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[68]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[69])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[70]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[71])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[72]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[73])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[74]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[75])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[76]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[77])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[78]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[79])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[80]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[81])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[82]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[83])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[84]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[85])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[86]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[87])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[88]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[89])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[90]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[91])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[92]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[93])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[94]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[95])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[96]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[97])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[98]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[99])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[100]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[101])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[102]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[103])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[104]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[105])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[106]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[107])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[108]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[109])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[110]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[111])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[112]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[113])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[114]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[115])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[116]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[117])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[118]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[119])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[120]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[121])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[122]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[123])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[124]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[125])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[126]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[127])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[128]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[129])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[130]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[131])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[132]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[133])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[134]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[135])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[136]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[137])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[138]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[139])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[140]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[141])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[142]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[143])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[144]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[145])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[146]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[147])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[148]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[149])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[150]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[151])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[152]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[153])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[154]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[155])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[156]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[157])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[158]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[159])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[160]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[161])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[162]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[163])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[164]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[165])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[166]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[167])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[168]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[169])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[170]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[171])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[172]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[173])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[174]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[175])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[176]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[177])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[178]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[179])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[180]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[181])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[182]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[183])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[184]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[185])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[186]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[187])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[188]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[189])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[190]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[191])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[192]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[193])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[194]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[195])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[196]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[197])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[198]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[199])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[200]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[201])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[202]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[203])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[204]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[205])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[206]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[207])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[208]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[209])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[210]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[211])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[212]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[213])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[214]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[215])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[216]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[217])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[218]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[219])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[220]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[221])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[222]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[223])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[224]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[225])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[226]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[227])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[228]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[229])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[230]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[231])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[232]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[233])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[234]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[235])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[236]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[237])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[238]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[239])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[240]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[241])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[242]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[243])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[244]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[245])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[246]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[247])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[248]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[249])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[250]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[251])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[252]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[253])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[254]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[255])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[256]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[257])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[258]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[259])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[260]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[261])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[262]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[263])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[264]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[265])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[266]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[267])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[268]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[269])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[270]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[271])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[272]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[273])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[274]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[275])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[276]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[277])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[278]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[279])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[280]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[281])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[282]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[283])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[284]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[285])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[286]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[287])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[288]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[289])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[290]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[291])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[292]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[293])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[294]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[295])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[296]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[297])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[298]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[299])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[300]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[301])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[302]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[303])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[304]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[305])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[306]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[307])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[308]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[309])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[310]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[311])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[312]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[313])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[314]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[315])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[316]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[317])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[318]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[319])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[320]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[321])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[322]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[323])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[324]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[325])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[326]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[327])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[328]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[329])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[330]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[331])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[332]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[333])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[334]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[335])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[336]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[337])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[338]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[339])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[340]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[341])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[342]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[343])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[344]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[345])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[346]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[347])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[348]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[349])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[350]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[351])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[352]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[353])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[354]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[355])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[356]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[357])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[358]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[359])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[360]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[361])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[362]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[363])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[364]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[365])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[366]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[367])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[368]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[369])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[370]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[371])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[372]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[373])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[374]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[375])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[376]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[377])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[378]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[379])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[380]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[381])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[382]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[383])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[384]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[385])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[386]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[387])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[388]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[389])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[390]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[391])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[392]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[393])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[394]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[395])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[396]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[397])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[398]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[399])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[400]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[401])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[402]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[403])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[404]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[405])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[406]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[407])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[408]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[409])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[410]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[411])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[412]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[413])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[414]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[415])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[416]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[417])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[418]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[419])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[420]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[421])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[422]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[423])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[424]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[425])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[426]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[427])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[428]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[429])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[430]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[431])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[432]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[433])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[434]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[435])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[436]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[437])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[438]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[439])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[440]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[441])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[442]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[443])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[444]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[445])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[446]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[447])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[448]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[449])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[450]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[451])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[452]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[453])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[454]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[455])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[456]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[457])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[458]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[459])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[460]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[461])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[462]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[463])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[464]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[465])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[466]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[467])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[468]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[469])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[470]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[471])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[472]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[473])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[474]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[475])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[476]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[477])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[478]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[479])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[480]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[481])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[482]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[483])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[484]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[485])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[486]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[487])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[488]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[489])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[490]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[491])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[492]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[493])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[494]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[495])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[496]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[497])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[498]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[499])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[500]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[501])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[502]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[503])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[504]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[505])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[506]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[507])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[508]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[509])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[510]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[511])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[512]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[513])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[514]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[515])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[516]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[517])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[518]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[519])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[520]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[521])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[522]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[523])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[524]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[525])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[526]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[527])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[528]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[529])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[530]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[531])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[532]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[533])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[534]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[535])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[536]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[537])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[538]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[539])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[540]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[541])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[542]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[543])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[544]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[545])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[546]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[547])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[548]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[549])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[550]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[551])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[552]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[553])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[554]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[555])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[556]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[557])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[558]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[559])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[560]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[561])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[562]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[563])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[564]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[565])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[566]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[567])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[568]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[569])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[570]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[571])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[572]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[573])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[574]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[575])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[576]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[577])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[578]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[579])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[580]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[581])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[582]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[583])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[584]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[585])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[586]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[587])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[588]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[589])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[590]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[591])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[592]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[593])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[594]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[595])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[596]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[597])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[598]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[599])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[600]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[601])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[602]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[603])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[604]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[605])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[606]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[607])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[608]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[609])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[610]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[611])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[612]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[613])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[614]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[615])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[616]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[617])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[618]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[619])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[620]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[621])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[622]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[623])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[624]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[625])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[626]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[627])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[628]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[629])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[630]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[631])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[632]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[633])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[634]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[635])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[636]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[637])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[638]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[639])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[640]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[641])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[642]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[643])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[644]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[645])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[646]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[647])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[648]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[649])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[650]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[651])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[652]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[653])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[654]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[655])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[656]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[657])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[658]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[659])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[660]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[661])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[662]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[663])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[664]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[665])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[666]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[667])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[668]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[669])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[670]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[671])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[672]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[673])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[674]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[675])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[676]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[677])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[678]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[679])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[680]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[681])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[682]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[683])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[684]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[685])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[686]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[687])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[688]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[689])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[690]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[691])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[692]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[693])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[694]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[695])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[696]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[697])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[698]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[699])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[700]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[701])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[702]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[703])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[704]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[705])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[706]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[707])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[708]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[709])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[710]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[711])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[712]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[713])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[714]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[715])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[716]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[717])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[718]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[719])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[720]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[721])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[722]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[723])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[724]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[725])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[726]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[727])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[728]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[729])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[730]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[731])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[732]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[733])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[734]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[735])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[736]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[737])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[738]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[739])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[740]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[741])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[742]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[743])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[744]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[745])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[746]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[747])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[748]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[749])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[750]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[751])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[752]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[753])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[754]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[755])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[756]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[757])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[758]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[759])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[760]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[761])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[762]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[763])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[764]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[765])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[766]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[767])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[768]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[769])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[770]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[771])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[772]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[773])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[774]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[775])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[776]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[777])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[778]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[779])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[780]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[781])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[782]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[783])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[784]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[785])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[786]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[787])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[788]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[789])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[790]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[791])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[792]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[793])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[794]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[795])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[796]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[797])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[798]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[799])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[800]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[801])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[802]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[803])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[804]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[805])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[806]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[807])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[808]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[809])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[810]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[811])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[812]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[813])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[814]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[815])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[816]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[817])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[818]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[819])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[820]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[821])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[822]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[823])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[824]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[825])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[826]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[827])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[828]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[829])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[830]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[831])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[832]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[833])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[834]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[835])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[836]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[837])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[838]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[839])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[840]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[841])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[842]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[843])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[844]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[845])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[846]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[847])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[848]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[849])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[850]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[851])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[852]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[853])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[854]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[855])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[856]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[857])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[858]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[859])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[860]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[861])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[862]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[863])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[864]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[865])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[866]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[867])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[868]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[869])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[870]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[871])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[872]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[873])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[874]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[875])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[876]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[877])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[878]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[879])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[880]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[881])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[882]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[883])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[884]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[885])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[886]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[887])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[888]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[889])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[890]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[891])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[892]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[893])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[894]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[895])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[896]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[897])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[898]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[899])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[900]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[901])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[902]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[903])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[904]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[905])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[906]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[907])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[908]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[909])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[910]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[911])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[912]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[913])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[914]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[915])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[916]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[917])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[918]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[919])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[920]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[921])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[922]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[923])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[924]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[925])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[926]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[927])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[928]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[929])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[930]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[931])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[932]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[933])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[934]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[935])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[936]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[937])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[938]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[939])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[940]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[941])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[942]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[943])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[944]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[945])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[946]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[947])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[948]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[949])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[950]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[951])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[952]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[953])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[954]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[955])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[956]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[957])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[958]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[959])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[960]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[961])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[962]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[963])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[964]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[965])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[966]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[967])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[968]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[969])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[970]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[971])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[972]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[973])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[974]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[975])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[976]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[977])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[978]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[979])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[980]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[981])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[982]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[983])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[984]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[985])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[986]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[987])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[988]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[989])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[990]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[991])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[992]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[993])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[994]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[995])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[996]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[997])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[998]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[999])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1000]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1001])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1002]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1003])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1004]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1005])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1006]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1007])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1008]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1009])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1010]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1011])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1012]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1013])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1014]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1015])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1016]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1017])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1018]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1019])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1020]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1021])
      | (~ (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1086])));
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva = conv_s2s_64_65(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1086:1023])
      + conv_u2s_1_65(mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_and_nl);
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva = nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[64:0];
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1022])
      & ((IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[0]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[2]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[3])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[4]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[5])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[6]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[7])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[8]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[9])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[10]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[11])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[12]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[13])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[14]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[15])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[16]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[17])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[18]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[19])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[20]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[21])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[22]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[23])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[24]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[25])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[26]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[27])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[28]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[29])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[30]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[31])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[32]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[33])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[34]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[35])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[36]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[37])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[38]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[39])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[40]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[41])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[42]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[43])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[44]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[45])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[46]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[47])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[48]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[49])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[50]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[51])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[52]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[53])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[54]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[55])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[56]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[57])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[58]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[59])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[60]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[61])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[62]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[63])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[64]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[65])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[66]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[67])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[68]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[69])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[70]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[71])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[72]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[73])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[74]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[75])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[76]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[77])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[78]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[79])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[80]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[81])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[82]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[83])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[84]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[85])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[86]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[87])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[88]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[89])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[90]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[91])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[92]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[93])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[94]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[95])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[96]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[97])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[98]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[99])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[100]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[101])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[102]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[103])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[104]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[105])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[106]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[107])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[108]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[109])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[110]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[111])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[112]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[113])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[114]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[115])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[116]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[117])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[118]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[119])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[120]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[121])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[122]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[123])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[124]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[125])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[126]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[127])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[128]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[129])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[130]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[131])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[132]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[133])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[134]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[135])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[136]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[137])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[138]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[139])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[140]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[141])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[142]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[143])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[144]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[145])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[146]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[147])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[148]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[149])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[150]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[151])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[152]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[153])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[154]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[155])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[156]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[157])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[158]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[159])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[160]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[161])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[162]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[163])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[164]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[165])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[166]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[167])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[168]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[169])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[170]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[171])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[172]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[173])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[174]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[175])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[176]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[177])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[178]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[179])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[180]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[181])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[182]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[183])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[184]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[185])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[186]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[187])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[188]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[189])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[190]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[191])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[192]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[193])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[194]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[195])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[196]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[197])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[198]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[199])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[200]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[201])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[202]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[203])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[204]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[205])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[206]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[207])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[208]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[209])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[210]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[211])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[212]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[213])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[214]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[215])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[216]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[217])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[218]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[219])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[220]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[221])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[222]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[223])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[224]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[225])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[226]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[227])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[228]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[229])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[230]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[231])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[232]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[233])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[234]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[235])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[236]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[237])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[238]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[239])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[240]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[241])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[242]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[243])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[244]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[245])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[246]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[247])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[248]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[249])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[250]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[251])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[252]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[253])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[254]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[255])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[256]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[257])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[258]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[259])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[260]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[261])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[262]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[263])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[264]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[265])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[266]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[267])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[268]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[269])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[270]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[271])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[272]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[273])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[274]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[275])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[276]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[277])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[278]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[279])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[280]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[281])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[282]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[283])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[284]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[285])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[286]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[287])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[288]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[289])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[290]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[291])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[292]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[293])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[294]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[295])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[296]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[297])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[298]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[299])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[300]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[301])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[302]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[303])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[304]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[305])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[306]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[307])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[308]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[309])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[310]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[311])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[312]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[313])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[314]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[315])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[316]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[317])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[318]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[319])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[320]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[321])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[322]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[323])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[324]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[325])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[326]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[327])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[328]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[329])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[330]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[331])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[332]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[333])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[334]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[335])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[336]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[337])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[338]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[339])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[340]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[341])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[342]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[343])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[344]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[345])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[346]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[347])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[348]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[349])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[350]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[351])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[352]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[353])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[354]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[355])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[356]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[357])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[358]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[359])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[360]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[361])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[362]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[363])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[364]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[365])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[366]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[367])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[368]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[369])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[370]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[371])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[372]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[373])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[374]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[375])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[376]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[377])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[378]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[379])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[380]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[381])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[382]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[383])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[384]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[385])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[386]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[387])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[388]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[389])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[390]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[391])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[392]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[393])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[394]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[395])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[396]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[397])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[398]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[399])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[400]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[401])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[402]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[403])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[404]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[405])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[406]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[407])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[408]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[409])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[410]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[411])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[412]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[413])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[414]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[415])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[416]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[417])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[418]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[419])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[420]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[421])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[422]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[423])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[424]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[425])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[426]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[427])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[428]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[429])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[430]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[431])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[432]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[433])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[434]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[435])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[436]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[437])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[438]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[439])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[440]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[441])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[442]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[443])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[444]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[445])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[446]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[447])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[448]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[449])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[450]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[451])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[452]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[453])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[454]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[455])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[456]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[457])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[458]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[459])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[460]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[461])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[462]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[463])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[464]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[465])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[466]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[467])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[468]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[469])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[470]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[471])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[472]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[473])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[474]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[475])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[476]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[477])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[478]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[479])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[480]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[481])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[482]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[483])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[484]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[485])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[486]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[487])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[488]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[489])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[490]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[491])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[492]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[493])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[494]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[495])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[496]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[497])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[498]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[499])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[500]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[501])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[502]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[503])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[504]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[505])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[506]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[507])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[508]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[509])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[510]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[511])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[512]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[513])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[514]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[515])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[516]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[517])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[518]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[519])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[520]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[521])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[522]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[523])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[524]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[525])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[526]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[527])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[528]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[529])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[530]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[531])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[532]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[533])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[534]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[535])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[536]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[537])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[538]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[539])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[540]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[541])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[542]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[543])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[544]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[545])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[546]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[547])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[548]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[549])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[550]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[551])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[552]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[553])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[554]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[555])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[556]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[557])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[558]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[559])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[560]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[561])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[562]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[563])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[564]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[565])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[566]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[567])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[568]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[569])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[570]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[571])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[572]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[573])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[574]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[575])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[576]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[577])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[578]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[579])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[580]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[581])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[582]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[583])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[584]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[585])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[586]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[587])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[588]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[589])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[590]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[591])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[592]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[593])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[594]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[595])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[596]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[597])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[598]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[599])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[600]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[601])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[602]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[603])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[604]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[605])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[606]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[607])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[608]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[609])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[610]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[611])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[612]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[613])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[614]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[615])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[616]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[617])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[618]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[619])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[620]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[621])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[622]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[623])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[624]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[625])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[626]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[627])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[628]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[629])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[630]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[631])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[632]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[633])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[634]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[635])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[636]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[637])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[638]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[639])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[640]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[641])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[642]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[643])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[644]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[645])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[646]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[647])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[648]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[649])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[650]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[651])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[652]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[653])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[654]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[655])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[656]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[657])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[658]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[659])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[660]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[661])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[662]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[663])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[664]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[665])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[666]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[667])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[668]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[669])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[670]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[671])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[672]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[673])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[674]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[675])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[676]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[677])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[678]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[679])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[680]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[681])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[682]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[683])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[684]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[685])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[686]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[687])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[688]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[689])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[690]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[691])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[692]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[693])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[694]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[695])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[696]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[697])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[698]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[699])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[700]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[701])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[702]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[703])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[704]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[705])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[706]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[707])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[708]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[709])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[710]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[711])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[712]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[713])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[714]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[715])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[716]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[717])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[718]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[719])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[720]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[721])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[722]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[723])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[724]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[725])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[726]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[727])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[728]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[729])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[730]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[731])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[732]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[733])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[734]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[735])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[736]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[737])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[738]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[739])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[740]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[741])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[742]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[743])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[744]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[745])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[746]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[747])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[748]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[749])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[750]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[751])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[752]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[753])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[754]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[755])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[756]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[757])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[758]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[759])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[760]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[761])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[762]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[763])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[764]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[765])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[766]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[767])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[768]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[769])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[770]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[771])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[772]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[773])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[774]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[775])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[776]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[777])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[778]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[779])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[780]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[781])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[782]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[783])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[784]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[785])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[786]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[787])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[788]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[789])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[790]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[791])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[792]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[793])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[794]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[795])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[796]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[797])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[798]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[799])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[800]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[801])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[802]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[803])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[804]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[805])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[806]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[807])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[808]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[809])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[810]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[811])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[812]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[813])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[814]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[815])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[816]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[817])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[818]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[819])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[820]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[821])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[822]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[823])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[824]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[825])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[826]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[827])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[828]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[829])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[830]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[831])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[832]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[833])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[834]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[835])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[836]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[837])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[838]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[839])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[840]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[841])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[842]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[843])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[844]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[845])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[846]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[847])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[848]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[849])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[850]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[851])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[852]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[853])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[854]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[855])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[856]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[857])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[858]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[859])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[860]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[861])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[862]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[863])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[864]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[865])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[866]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[867])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[868]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[869])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[870]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[871])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[872]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[873])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[874]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[875])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[876]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[877])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[878]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[879])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[880]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[881])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[882]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[883])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[884]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[885])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[886]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[887])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[888]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[889])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[890]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[891])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[892]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[893])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[894]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[895])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[896]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[897])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[898]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[899])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[900]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[901])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[902]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[903])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[904]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[905])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[906]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[907])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[908]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[909])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[910]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[911])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[912]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[913])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[914]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[915])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[916]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[917])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[918]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[919])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[920]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[921])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[922]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[923])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[924]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[925])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[926]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[927])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[928]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[929])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[930]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[931])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[932]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[933])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[934]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[935])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[936]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[937])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[938]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[939])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[940]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[941])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[942]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[943])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[944]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[945])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[946]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[947])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[948]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[949])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[950]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[951])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[952]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[953])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[954]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[955])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[956]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[957])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[958]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[959])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[960]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[961])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[962]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[963])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[964]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[965])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[966]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[967])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[968]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[969])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[970]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[971])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[972]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[973])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[974]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[975])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[976]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[977])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[978]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[979])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[980]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[981])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[982]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[983])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[984]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[985])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[986]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[987])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[988]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[989])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[990]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[991])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[992]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[993])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[994]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[995])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[996]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[997])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[998]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[999])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1000]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1001])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1002]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1003])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1004]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1005])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1006]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1007])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1008]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1009])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1010]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1011])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1012]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1013])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1014]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1015])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1016]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1017])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1018]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1019])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1020]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1021])
      | (~ (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1086])));
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva = conv_s2s_64_65(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1086:1023])
      + conv_u2s_1_65(mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_and_nl);
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva = nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[64:0];
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1022])
      & ((IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[0]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[2]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[3])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[4]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[5])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[6]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[7])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[8]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[9])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[10]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[11])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[12]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[13])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[14]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[15])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[16]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[17])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[18]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[19])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[20]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[21])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[22]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[23])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[24]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[25])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[26]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[27])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[28]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[29])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[30]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[31])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[32]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[33])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[34]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[35])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[36]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[37])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[38]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[39])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[40]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[41])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[42]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[43])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[44]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[45])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[46]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[47])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[48]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[49])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[50]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[51])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[52]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[53])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[54]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[55])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[56]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[57])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[58]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[59])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[60]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[61])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[62]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[63])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[64]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[65])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[66]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[67])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[68]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[69])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[70]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[71])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[72]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[73])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[74]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[75])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[76]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[77])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[78]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[79])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[80]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[81])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[82]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[83])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[84]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[85])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[86]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[87])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[88]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[89])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[90]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[91])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[92]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[93])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[94]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[95])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[96]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[97])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[98]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[99])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[100]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[101])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[102]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[103])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[104]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[105])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[106]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[107])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[108]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[109])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[110]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[111])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[112]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[113])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[114]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[115])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[116]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[117])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[118]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[119])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[120]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[121])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[122]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[123])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[124]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[125])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[126]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[127])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[128]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[129])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[130]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[131])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[132]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[133])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[134]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[135])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[136]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[137])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[138]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[139])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[140]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[141])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[142]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[143])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[144]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[145])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[146]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[147])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[148]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[149])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[150]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[151])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[152]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[153])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[154]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[155])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[156]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[157])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[158]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[159])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[160]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[161])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[162]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[163])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[164]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[165])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[166]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[167])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[168]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[169])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[170]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[171])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[172]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[173])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[174]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[175])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[176]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[177])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[178]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[179])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[180]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[181])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[182]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[183])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[184]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[185])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[186]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[187])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[188]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[189])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[190]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[191])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[192]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[193])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[194]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[195])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[196]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[197])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[198]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[199])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[200]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[201])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[202]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[203])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[204]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[205])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[206]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[207])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[208]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[209])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[210]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[211])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[212]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[213])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[214]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[215])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[216]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[217])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[218]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[219])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[220]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[221])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[222]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[223])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[224]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[225])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[226]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[227])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[228]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[229])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[230]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[231])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[232]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[233])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[234]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[235])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[236]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[237])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[238]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[239])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[240]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[241])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[242]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[243])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[244]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[245])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[246]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[247])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[248]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[249])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[250]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[251])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[252]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[253])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[254]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[255])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[256]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[257])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[258]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[259])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[260]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[261])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[262]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[263])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[264]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[265])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[266]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[267])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[268]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[269])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[270]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[271])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[272]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[273])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[274]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[275])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[276]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[277])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[278]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[279])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[280]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[281])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[282]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[283])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[284]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[285])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[286]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[287])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[288]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[289])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[290]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[291])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[292]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[293])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[294]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[295])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[296]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[297])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[298]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[299])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[300]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[301])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[302]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[303])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[304]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[305])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[306]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[307])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[308]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[309])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[310]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[311])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[312]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[313])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[314]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[315])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[316]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[317])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[318]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[319])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[320]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[321])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[322]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[323])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[324]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[325])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[326]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[327])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[328]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[329])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[330]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[331])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[332]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[333])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[334]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[335])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[336]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[337])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[338]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[339])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[340]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[341])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[342]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[343])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[344]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[345])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[346]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[347])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[348]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[349])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[350]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[351])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[352]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[353])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[354]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[355])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[356]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[357])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[358]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[359])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[360]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[361])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[362]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[363])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[364]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[365])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[366]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[367])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[368]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[369])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[370]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[371])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[372]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[373])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[374]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[375])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[376]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[377])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[378]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[379])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[380]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[381])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[382]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[383])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[384]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[385])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[386]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[387])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[388]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[389])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[390]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[391])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[392]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[393])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[394]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[395])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[396]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[397])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[398]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[399])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[400]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[401])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[402]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[403])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[404]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[405])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[406]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[407])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[408]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[409])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[410]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[411])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[412]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[413])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[414]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[415])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[416]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[417])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[418]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[419])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[420]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[421])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[422]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[423])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[424]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[425])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[426]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[427])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[428]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[429])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[430]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[431])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[432]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[433])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[434]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[435])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[436]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[437])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[438]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[439])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[440]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[441])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[442]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[443])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[444]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[445])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[446]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[447])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[448]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[449])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[450]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[451])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[452]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[453])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[454]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[455])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[456]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[457])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[458]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[459])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[460]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[461])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[462]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[463])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[464]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[465])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[466]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[467])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[468]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[469])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[470]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[471])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[472]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[473])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[474]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[475])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[476]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[477])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[478]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[479])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[480]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[481])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[482]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[483])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[484]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[485])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[486]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[487])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[488]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[489])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[490]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[491])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[492]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[493])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[494]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[495])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[496]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[497])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[498]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[499])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[500]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[501])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[502]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[503])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[504]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[505])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[506]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[507])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[508]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[509])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[510]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[511])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[512]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[513])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[514]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[515])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[516]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[517])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[518]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[519])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[520]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[521])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[522]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[523])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[524]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[525])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[526]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[527])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[528]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[529])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[530]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[531])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[532]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[533])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[534]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[535])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[536]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[537])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[538]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[539])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[540]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[541])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[542]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[543])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[544]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[545])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[546]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[547])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[548]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[549])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[550]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[551])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[552]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[553])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[554]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[555])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[556]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[557])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[558]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[559])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[560]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[561])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[562]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[563])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[564]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[565])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[566]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[567])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[568]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[569])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[570]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[571])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[572]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[573])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[574]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[575])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[576]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[577])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[578]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[579])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[580]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[581])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[582]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[583])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[584]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[585])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[586]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[587])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[588]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[589])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[590]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[591])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[592]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[593])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[594]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[595])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[596]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[597])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[598]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[599])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[600]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[601])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[602]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[603])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[604]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[605])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[606]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[607])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[608]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[609])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[610]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[611])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[612]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[613])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[614]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[615])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[616]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[617])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[618]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[619])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[620]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[621])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[622]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[623])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[624]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[625])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[626]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[627])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[628]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[629])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[630]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[631])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[632]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[633])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[634]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[635])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[636]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[637])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[638]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[639])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[640]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[641])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[642]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[643])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[644]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[645])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[646]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[647])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[648]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[649])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[650]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[651])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[652]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[653])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[654]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[655])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[656]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[657])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[658]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[659])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[660]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[661])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[662]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[663])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[664]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[665])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[666]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[667])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[668]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[669])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[670]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[671])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[672]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[673])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[674]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[675])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[676]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[677])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[678]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[679])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[680]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[681])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[682]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[683])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[684]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[685])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[686]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[687])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[688]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[689])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[690]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[691])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[692]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[693])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[694]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[695])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[696]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[697])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[698]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[699])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[700]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[701])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[702]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[703])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[704]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[705])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[706]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[707])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[708]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[709])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[710]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[711])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[712]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[713])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[714]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[715])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[716]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[717])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[718]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[719])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[720]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[721])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[722]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[723])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[724]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[725])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[726]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[727])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[728]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[729])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[730]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[731])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[732]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[733])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[734]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[735])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[736]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[737])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[738]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[739])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[740]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[741])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[742]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[743])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[744]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[745])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[746]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[747])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[748]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[749])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[750]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[751])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[752]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[753])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[754]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[755])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[756]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[757])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[758]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[759])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[760]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[761])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[762]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[763])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[764]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[765])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[766]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[767])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[768]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[769])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[770]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[771])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[772]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[773])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[774]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[775])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[776]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[777])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[778]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[779])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[780]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[781])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[782]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[783])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[784]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[785])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[786]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[787])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[788]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[789])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[790]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[791])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[792]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[793])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[794]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[795])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[796]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[797])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[798]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[799])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[800]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[801])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[802]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[803])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[804]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[805])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[806]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[807])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[808]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[809])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[810]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[811])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[812]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[813])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[814]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[815])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[816]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[817])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[818]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[819])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[820]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[821])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[822]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[823])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[824]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[825])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[826]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[827])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[828]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[829])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[830]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[831])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[832]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[833])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[834]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[835])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[836]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[837])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[838]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[839])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[840]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[841])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[842]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[843])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[844]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[845])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[846]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[847])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[848]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[849])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[850]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[851])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[852]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[853])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[854]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[855])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[856]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[857])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[858]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[859])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[860]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[861])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[862]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[863])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[864]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[865])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[866]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[867])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[868]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[869])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[870]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[871])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[872]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[873])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[874]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[875])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[876]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[877])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[878]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[879])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[880]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[881])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[882]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[883])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[884]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[885])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[886]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[887])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[888]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[889])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[890]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[891])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[892]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[893])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[894]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[895])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[896]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[897])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[898]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[899])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[900]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[901])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[902]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[903])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[904]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[905])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[906]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[907])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[908]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[909])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[910]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[911])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[912]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[913])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[914]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[915])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[916]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[917])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[918]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[919])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[920]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[921])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[922]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[923])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[924]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[925])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[926]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[927])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[928]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[929])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[930]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[931])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[932]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[933])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[934]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[935])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[936]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[937])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[938]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[939])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[940]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[941])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[942]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[943])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[944]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[945])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[946]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[947])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[948]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[949])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[950]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[951])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[952]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[953])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[954]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[955])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[956]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[957])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[958]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[959])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[960]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[961])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[962]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[963])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[964]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[965])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[966]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[967])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[968]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[969])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[970]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[971])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[972]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[973])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[974]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[975])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[976]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[977])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[978]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[979])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[980]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[981])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[982]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[983])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[984]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[985])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[986]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[987])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[988]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[989])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[990]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[991])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[992]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[993])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[994]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[995])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[996]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[997])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[998]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[999])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1000]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1001])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1002]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1003])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1004]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1005])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1006]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1007])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1008]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1009])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1010]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1011])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1012]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1013])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1014]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1015])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1016]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1017])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1018]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1019])
      | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1020]) | (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1021])
      | (~ (IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1086])));
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva = conv_s2s_64_65(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1086:1023])
      + conv_u2s_1_65(mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_and_nl);
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva = nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[64:0];
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_1_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = readslicef_8_1_7((mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_743_nl = (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign mux_233_nl = MUX_s_1_2_2((mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_1_sva[47]), or_743_nl);
  assign FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_1_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_1_sva_mx1[46:1]), mux_233_nl);
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_2_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = readslicef_8_1_7((mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_744_nl = (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign mux_234_nl = MUX_s_1_2_2((mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_2_sva[47]), or_744_nl);
  assign FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_2_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_2_sva_mx1[46:1]), mux_234_nl);
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_3_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = readslicef_8_1_7((mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign or_745_nl = (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign mux_235_nl = MUX_s_1_2_2((mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_3_sva[47]), or_745_nl);
  assign FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_3_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_3_sva_mx1[46:1]), mux_235_nl);
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_8U_23U_p_expo_sva_1_mx0w0[7:1])})
      + 8'b1;
  assign mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0];
  assign mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = readslicef_8_1_7((mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl));
  assign mux_236_nl = MUX_s_1_2_2((mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
      (FpMul_8U_23U_p_mant_p1_sva[47]), or_430_cse);
  assign FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0 = MUX_v_46_2_2((FpMul_8U_23U_p_mant_p1_sva_mx1[45:0]),
      (FpMul_8U_23U_p_mant_p1_sva_mx1[46:1]), mux_236_nl);
  assign asn_156 = mul_mul_else_unequal_tmp_1 & (~ mul_mul_land_lpi_1_dfm_6) & (~
      io_read_cfg_mul_bypass_rsc_svs_5);
  assign asn_158 = mul_mul_land_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5;
  assign asn_160 = mul_mul_else_unequal_tmp_1 & (~ mul_mul_land_1_lpi_1_dfm_6) &
      (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign asn_162 = mul_mul_land_1_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5;
  assign asn_164 = mul_mul_else_unequal_tmp_1 & (~ mul_mul_land_3_lpi_1_dfm_6) &
      (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign asn_166 = mul_mul_land_3_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5;
  assign asn_168 = mul_mul_else_unequal_tmp_1 & (~ mul_mul_land_2_lpi_1_dfm_6) &
      (~ io_read_cfg_mul_bypass_rsc_svs_5);
  assign asn_170 = mul_mul_land_2_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5;
  assign and_18_tmp = main_stage_v_1 & or_11_cse & or_12_cse & or_13_cse & or_14_cse
      & or_15_cse & or_16_cse & or_74_cse;
  assign else_mux_3_tmp_30_23 = MUX_v_8_2_2((cfg_mul_op_1_sva_1[30:23]), (chn_mul_op_rsci_d_mxwt[126:119]),
      cfg_mul_src_1_sva_1);
  assign else_mux_2_tmp_30_23 = MUX_v_8_2_2((cfg_mul_op_1_sva_1[30:23]), (chn_mul_op_rsci_d_mxwt[94:87]),
      cfg_mul_src_1_sva_1);
  assign else_mux_1_tmp_30_23 = MUX_v_8_2_2((cfg_mul_op_1_sva_1[30:23]), (chn_mul_op_rsci_d_mxwt[62:55]),
      cfg_mul_src_1_sva_1);
  assign else_mux_tmp_30_23 = MUX_v_8_2_2((cfg_mul_op_1_sva_1[30:23]), (chn_mul_op_rsci_d_mxwt[30:23]),
      cfg_mul_src_1_sva_1);
  assign or_tmp_1 = io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_1_lpi_1_dfm_st_1;
  assign or_19_nl = mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_land_1_lpi_1_dfm_4
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp | (~ mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign mux_5_nl = MUX_s_1_2_2(or_469_cse, (or_19_nl), nor_20_cse);
  assign nor_nl = ~(or_tmp_1 | (mux_5_nl));
  assign nor_331_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt);
  assign not_tmp_2 = MUX_s_1_2_2((nor_331_nl), (nor_nl), and_18_tmp);
  assign or_26_nl = mul_mul_land_1_lpi_1_dfm_st_4 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2);
  assign mux_7_itm = MUX_s_1_2_2((or_26_nl), or_tmp_1, and_18_tmp);
  assign or_tmp_12 = mul_mul_land_1_lpi_1_dfm_st_1 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | IsZero_8U_23U_land_1_lpi_1_dfm_4 | mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  assign or_tmp_15 = io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_2_lpi_1_dfm_st_1;
  assign or_34_nl = mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_land_2_lpi_1_dfm_4
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp | (~ mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign mux_10_nl = MUX_s_1_2_2(or_482_cse, (or_34_nl), nor_20_cse);
  assign nor_326_nl = ~(or_tmp_15 | (mux_10_nl));
  assign nor_327_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt);
  assign not_tmp_8 = MUX_s_1_2_2((nor_327_nl), (nor_326_nl), and_18_tmp);
  assign or_40_nl = mul_mul_land_2_lpi_1_dfm_st_4 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2);
  assign mux_12_itm = MUX_s_1_2_2((or_40_nl), or_tmp_15, and_18_tmp);
  assign or_tmp_26 = mul_mul_land_2_lpi_1_dfm_st_1 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | IsZero_8U_23U_land_2_lpi_1_dfm_4 | mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  assign or_tmp_29 = io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_3_lpi_1_dfm_st_1;
  assign or_48_nl = mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_land_3_lpi_1_dfm_4
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp | (~ mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign mux_15_nl = MUX_s_1_2_2(or_490_cse, (or_48_nl), nor_20_cse);
  assign nor_324_nl = ~(or_tmp_29 | (mux_15_nl));
  assign nor_325_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt);
  assign not_tmp_12 = MUX_s_1_2_2((nor_325_nl), (nor_324_nl), and_18_tmp);
  assign or_54_nl = mul_mul_land_3_lpi_1_dfm_st_4 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2);
  assign mux_17_itm = MUX_s_1_2_2((or_54_nl), or_tmp_29, and_18_tmp);
  assign or_tmp_40 = mul_mul_land_3_lpi_1_dfm_st_1 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | IsZero_8U_23U_land_3_lpi_1_dfm_4 | mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  assign nor_321_nl = ~(mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_land_lpi_1_dfm_4
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp | (~ mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1)
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_lpi_1_dfm_st_1);
  assign nor_322_nl = ~((~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_lpi_1_dfm_st_1);
  assign mux_20_nl = MUX_s_1_2_2((nor_322_nl), (nor_321_nl), nor_20_cse);
  assign nor_323_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt);
  assign not_tmp_15 = MUX_s_1_2_2((nor_323_nl), (mux_20_nl), and_18_tmp);
  assign or_tmp_46 = mul_mul_land_lpi_1_dfm_st_1 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_65_nl = (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mul_mul_land_lpi_1_dfm_st_4 | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2);
  assign mux_22_itm = MUX_s_1_2_2((or_65_nl), or_tmp_46, and_18_tmp);
  assign or_tmp_51 = mul_mul_land_lpi_1_dfm_st_1 | io_read_cfg_mul_bypass_rsc_svs_st_1
      | mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp
      | IsZero_8U_23U_land_lpi_1_dfm_4;
  assign or_tmp_59 = io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4;
  assign or_tmp_75 = io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4;
  assign or_tmp_91 = io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4;
  assign or_tmp_107 = io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4;
  assign or_tmp_123 = io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5;
  assign or_tmp_128 = FpMul_8U_23U_FpMul_8U_23U_and_itm | FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign or_tmp_132 = (mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2
      & FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3)
      | FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2;
  assign or_tmp_133 = FpMul_8U_23U_lor_6_lpi_1_dfm_7 | FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  assign or_tmp_146 = io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5;
  assign or_tmp_167 = nor_143_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2);
  assign or_tmp_173 = io_read_cfg_mul_bypass_rsc_svs_5 | (~ main_stage_v_3);
  assign or_189_cse = io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2);
  assign mux_tmp_46 = MUX_s_1_2_2(or_tmp_173, or_189_cse, or_74_cse);
  assign or_187_nl = mul_mul_land_1_lpi_1_dfm_st_5 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_5 | (~ main_stage_v_3);
  assign mux_52_nl = MUX_s_1_2_2(mux_tmp_46, or_tmp_167, mul_mul_land_1_lpi_1_dfm_st_5);
  assign mux_tmp_48 = MUX_s_1_2_2((mux_52_nl), (or_187_nl), mul_mul_land_1_lpi_1_dfm_st_4);
  assign nor_285_nl = ~(mul_mul_land_1_lpi_1_dfm_6 | mul_mul_land_1_lpi_1_dfm_st_5
      | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3));
  assign nor_286_nl = ~(nor_143_cse | mul_mul_land_1_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2));
  assign nor_288_nl = ~(mul_mul_land_1_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2));
  assign nor_289_nl = ~(io_read_cfg_mul_bypass_rsc_svs_5 | (~ main_stage_v_3));
  assign mux_56_nl = MUX_s_1_2_2((nor_289_nl), (nor_288_nl), or_74_cse);
  assign or_193_nl = mul_mul_land_1_lpi_1_dfm_6 | mul_mul_land_1_lpi_1_dfm_st_5;
  assign mux_57_nl = MUX_s_1_2_2((mux_56_nl), (nor_286_nl), or_193_nl);
  assign not_tmp_54 = MUX_s_1_2_2((mux_57_nl), (nor_285_nl), mul_mul_land_1_lpi_1_dfm_st_4);
  assign nor_283_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5);
  assign nor_284_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_8 | mul_mul_land_1_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_7);
  assign not_tmp_55 = MUX_s_1_2_2((nor_284_nl), (nor_283_nl), or_74_cse);
  assign or_tmp_211 = FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign or_tmp_216 = FpMul_8U_23U_FpMul_8U_23U_and_12_itm | FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign or_tmp_235 = io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign or_tmp_252 = FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | mul_mul_land_2_lpi_1_dfm_st_4;
  assign or_tmp_256 = mul_mul_land_2_lpi_1_dfm_st_5 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_5 | (~ main_stage_v_3);
  assign mux_tmp_78 = MUX_s_1_2_2(mux_tmp_46, or_tmp_167, mul_mul_land_2_lpi_1_dfm_st_5);
  assign nor_248_nl = ~(mul_mul_land_2_lpi_1_dfm_st_5 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | mul_mul_land_2_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3));
  assign nor_249_nl = ~(nor_143_cse | mul_mul_land_2_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2));
  assign nor_251_nl = ~(mul_mul_land_2_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2));
  assign nor_252_nl = ~(mul_mul_land_2_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3));
  assign mux_86_nl = MUX_s_1_2_2((nor_252_nl), (nor_251_nl), or_74_cse);
  assign mux_87_nl = MUX_s_1_2_2((mux_86_nl), (nor_249_nl), mul_mul_land_2_lpi_1_dfm_st_5);
  assign not_tmp_81 = MUX_s_1_2_2((mux_87_nl), (nor_248_nl), mul_mul_land_2_lpi_1_dfm_st_4);
  assign nor_246_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_7
      | mul_mul_land_2_lpi_1_dfm_5);
  assign nor_247_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_8 | mul_mul_land_2_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_7);
  assign not_tmp_82 = MUX_s_1_2_2((nor_247_nl), (nor_246_nl), or_74_cse);
  assign mux_94_itm = MUX_s_1_2_2(mux_tmp_78, or_tmp_256, mul_mul_land_2_lpi_1_dfm_st_4);
  assign or_tmp_291 = FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign or_tmp_296 = FpMul_8U_23U_FpMul_8U_23U_and_13_itm | FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign or_tmp_315 = io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign or_tmp_332 = FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | mul_mul_land_3_lpi_1_dfm_st_4;
  assign or_tmp_336 = mul_mul_land_3_lpi_1_dfm_st_5 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_5 | (~ main_stage_v_3);
  assign mux_tmp_109 = MUX_s_1_2_2(mux_tmp_46, or_tmp_167, mul_mul_land_3_lpi_1_dfm_st_5);
  assign nor_211_nl = ~(mul_mul_land_3_lpi_1_dfm_st_5 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | mul_mul_land_3_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3));
  assign nor_212_nl = ~(nor_143_cse | mul_mul_land_3_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2));
  assign nor_214_nl = ~(mul_mul_land_3_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2));
  assign nor_215_nl = ~(mul_mul_land_3_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3));
  assign mux_117_nl = MUX_s_1_2_2((nor_215_nl), (nor_214_nl), or_74_cse);
  assign mux_118_nl = MUX_s_1_2_2((mux_117_nl), (nor_212_nl), mul_mul_land_3_lpi_1_dfm_st_5);
  assign not_tmp_106 = MUX_s_1_2_2((mux_118_nl), (nor_211_nl), mul_mul_land_3_lpi_1_dfm_st_4);
  assign nor_209_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_7
      | mul_mul_land_3_lpi_1_dfm_5);
  assign nor_210_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_8 | mul_mul_land_3_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_7);
  assign not_tmp_107 = MUX_s_1_2_2((nor_210_nl), (nor_209_nl), or_74_cse);
  assign mux_125_itm = MUX_s_1_2_2(mux_tmp_109, or_tmp_336, mul_mul_land_3_lpi_1_dfm_st_4);
  assign or_tmp_371 = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign or_tmp_376 = FpMul_8U_23U_FpMul_8U_23U_and_14_itm | FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign not_tmp_121 = ~(mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
      & main_stage_v_2);
  assign or_tmp_395 = io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_1_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign or_tmp_411 = nor_143_cse | mul_mul_land_lpi_1_dfm_st_4 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2);
  assign or_tmp_415 = mul_mul_land_lpi_1_dfm_st_5 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_5 | (~ main_stage_v_3);
  assign or_435_nl = or_tmp_107 | (~ main_stage_v_2);
  assign mux_144_nl = MUX_s_1_2_2(or_tmp_173, (or_435_nl), or_74_cse);
  assign mux_tmp_140 = MUX_s_1_2_2((mux_144_nl), or_tmp_411, mul_mul_land_lpi_1_dfm_st_5);
  assign nor_177_nl = ~(nor_143_cse | mul_mul_land_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_lpi_1_dfm_st_4 | (~ main_stage_v_2));
  assign nor_179_nl = ~(mul_mul_land_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_lpi_1_dfm_st_4 | (~ main_stage_v_2));
  assign nor_180_nl = ~(mul_mul_land_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3));
  assign mux_150_nl = MUX_s_1_2_2((nor_180_nl), (nor_179_nl), or_74_cse);
  assign not_tmp_129 = MUX_s_1_2_2((mux_150_nl), (nor_177_nl), mul_mul_land_lpi_1_dfm_st_5);
  assign nor_175_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | IsNaN_8U_23U_1_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_7
      | mul_mul_land_lpi_1_dfm_5);
  assign nor_176_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_8 | mul_mul_land_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_lpi_1_dfm_7);
  assign not_tmp_130 = MUX_s_1_2_2((nor_176_nl), (nor_175_nl), or_74_cse);
  assign or_tmp_461 = (~((chn_mul_in_rsci_d_mxwt[95]) | (chn_mul_in_rsci_d_mxwt[31])
      | (chn_mul_in_rsci_d_mxwt[63]) | (chn_mul_in_rsci_d_mxwt[127]) | (~ cfg_mul_prelu_rsci_d)))
      | cfg_mul_bypass_rsci_d;
  assign and_dcpl_3 = and_20_tmp & (cfg_precision==2'b10);
  assign and_dcpl_4 = ~(mul_mul_land_1_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d);
  assign and_dcpl_6 = or_27_cse & and_20_tmp;
  assign and_dcpl_8 = ~(mul_mul_land_2_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d);
  assign and_dcpl_11 = ~(mul_mul_land_3_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d);
  assign and_dcpl_14 = ~(mul_mul_land_lpi_1_dfm_mx1w0 | cfg_mul_bypass_rsci_d);
  assign or_tmp_517 = FpMul_8U_23U_FpMul_8U_23U_and_14_itm | (~ or_tmp_411);
  assign and_tmp_5 = FpMul_8U_23U_FpMul_8U_23U_and_14_itm & or_tmp_411;
  assign and_dcpl_22 = main_stage_v_3 & (~ io_read_cfg_mul_bypass_rsc_svs_5) & or_74_cse;
  assign and_dcpl_23 = (~ chn_mul_out_rsci_bawt) & reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_24 = or_74_cse & main_stage_v_3;
  assign and_dcpl_26 = (~ main_stage_v_3) & chn_mul_out_rsci_bawt & reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_27 = (~ cfg_mul_bypass_rsci_d) & and_20_tmp;
  assign or_dcpl_8 = cfg_mul_bypass_rsci_d | (~ and_20_tmp);
  assign and_dcpl_30 = (~ io_read_cfg_mul_bypass_rsc_svs_st_1) & cfg_mul_src_1_sva_st_1
      & and_18_tmp;
  assign or_dcpl_13 = and_dcpl_23 | (~ main_stage_v_2);
  assign and_dcpl_37 = (cfg_precision==2'b10);
  assign and_dcpl_38 = and_dcpl_37 & and_18_tmp;
  assign and_dcpl_39 = or_27_cse & and_18_tmp;
  assign and_dcpl_45 = or_74_cse & (~ (cfg_precision[0]));
  assign and_dcpl_46 = and_dcpl_45 & (cfg_precision[1]) & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_6);
  assign and_dcpl_47 = or_74_cse & or_27_cse;
  assign and_dcpl_48 = and_dcpl_47 & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_6);
  assign and_dcpl_50 = and_dcpl_45 & (cfg_precision[1]) & IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign and_dcpl_51 = and_dcpl_47 & IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign and_dcpl_52 = or_74_cse & and_dcpl_37;
  assign and_dcpl_54 = and_dcpl_45 & (cfg_precision[1]) & (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_6);
  assign and_dcpl_55 = and_dcpl_47 & (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_6);
  assign and_dcpl_57 = and_dcpl_45 & (cfg_precision[1]) & IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign and_dcpl_58 = and_dcpl_47 & IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign and_dcpl_60 = and_dcpl_45 & (cfg_precision[1]) & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_6);
  assign and_dcpl_61 = and_dcpl_47 & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_6);
  assign and_dcpl_63 = and_dcpl_45 & (cfg_precision[1]) & IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign and_dcpl_64 = and_dcpl_47 & IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign and_dcpl_66 = and_dcpl_45 & (cfg_precision[1]) & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_6);
  assign and_dcpl_67 = and_dcpl_47 & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_6);
  assign and_dcpl_69 = and_dcpl_45 & (cfg_precision[1]) & IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign and_dcpl_70 = and_dcpl_47 & IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign or_dcpl_22 = or_dcpl_13 | or_tmp_59 | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3
      | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_27_cse;
  assign or_dcpl_23 = mul_mul_land_1_lpi_1_dfm_st_4 | (cfg_precision[0]);
  assign or_dcpl_26 = or_189_cse | and_dcpl_23;
  assign or_dcpl_27 = or_dcpl_26 | or_dcpl_23 | (~ (cfg_precision[1]));
  assign or_dcpl_37 = or_dcpl_13 | or_tmp_75 | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3
      | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_27_cse;
  assign or_dcpl_40 = or_dcpl_26 | mul_mul_land_2_lpi_1_dfm_st_4 | (cfg_precision!=2'b10);
  assign or_dcpl_50 = or_dcpl_13 | or_tmp_91 | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3
      | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_27_cse;
  assign or_dcpl_53 = or_dcpl_26 | mul_mul_land_3_lpi_1_dfm_st_4 | (cfg_precision!=2'b10);
  assign or_dcpl_63 = or_189_cse | mul_mul_land_lpi_1_dfm_st_4 | and_dcpl_23 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | or_27_cse;
  assign or_dcpl_66 = or_dcpl_26 | mul_mul_land_lpi_1_dfm_st_4 | (cfg_precision!=2'b10);
  assign or_dcpl_75 = IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp | mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  assign or_dcpl_81 = IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp | mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  assign or_dcpl_87 = IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp | mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  assign or_dcpl_93 = IsZero_8U_23U_land_lpi_1_dfm_4 | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign or_dcpl_96 = ~((cfg_precision[1]) & and_18_tmp);
  assign or_dcpl_99 = or_tmp_1 | (cfg_precision[0]) | or_dcpl_96;
  assign or_dcpl_102 = or_tmp_15 | (cfg_precision[0]) | or_dcpl_96;
  assign or_dcpl_105 = or_tmp_29 | (cfg_precision[0]) | or_dcpl_96;
  assign or_dcpl_108 = or_tmp_46 | (cfg_precision[0]) | or_dcpl_96;
  assign or_dcpl_110 = (~ and_20_tmp) | (cfg_precision!=2'b10);
  assign or_dcpl_125 = and_dcpl_37 | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign or_tmp_587 = and_20_tmp & (fsm_output[1]);
  assign or_tmp_588 = and_dcpl_27 & cfg_mul_src_rsci_d & (fsm_output[1]);
  assign or_tmp_591 = and_18_tmp & (fsm_output[1]);
  assign chn_mul_in_rsci_ld_core_psct_mx0c0 = and_20_tmp | (fsm_output[0]);
  assign chn_mul_op_rsci_ld_core_psct_mx0c1 = and_dcpl_30 & (or_dcpl_8 | (~ cfg_mul_src_rsci_d));
  assign main_stage_v_2_mx0c1 = or_74_cse & main_stage_v_2 & (~ and_18_tmp);
  assign main_stage_v_3_mx0c1 = main_stage_v_3 & (~ main_stage_v_2) & or_74_cse;
  assign main_stage_v_1_mx0c1 = (~ and_20_tmp) & and_18_tmp & (fsm_output[1]);
  assign cfg_mul_src_1_sva_st_1_mx0c1 = cfg_mul_bypass_rsci_d & and_20_tmp & (fsm_output[1]);
  assign chn_mul_in_rsci_oswt_unreg = or_tmp_587;
  assign chn_mul_op_rsci_oswt_unreg = and_dcpl_30;
  assign chn_mul_out_rsci_oswt_unreg = chn_mul_out_rsci_bawt & reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff = or_tmp_591;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_iswt0 <= 1'b0;
      reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      chn_mul_out_rsci_iswt0 <= 1'b0;
      chn_mul_op_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_mul_in_rsci_iswt0 <= ~((~ and_20_tmp) & (fsm_output[1]));
      reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse <= or_tmp_587;
      chn_mul_out_rsci_iswt0 <= and_dcpl_24;
      chn_mul_op_rsci_iswt0 <= or_tmp_588;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_mul_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_mul_in_rsci_ld_core_psct <= chn_mul_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_d_0 <= 1'b0;
      chn_mul_out_rsci_d_31 <= 1'b0;
      chn_mul_out_rsci_d_32 <= 1'b0;
      chn_mul_out_rsci_d_63 <= 1'b0;
      chn_mul_out_rsci_d_64 <= 1'b0;
      chn_mul_out_rsci_d_95 <= 1'b0;
      chn_mul_out_rsci_d_96 <= 1'b0;
      chn_mul_out_rsci_d_127 <= 1'b0;
    end
    else if ( chn_mul_out_and_cse ) begin
      chn_mul_out_rsci_d_0 <= MUX_s_1_2_2((MulIn_data_sva_133[0]), (mul_mul_mux_108_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_31 <= MUX_s_1_2_2((MulIn_data_sva_133[31]), (mul_mul_mux_109_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_32 <= MUX_s_1_2_2((MulIn_data_sva_133[32]), (mul_mul_mux_110_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_63 <= MUX_s_1_2_2((MulIn_data_sva_133[63]), (mul_mul_mux_111_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_64 <= MUX_s_1_2_2((MulIn_data_sva_133[64]), (mul_mul_mux_112_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_95 <= MUX_s_1_2_2((MulIn_data_sva_133[95]), (mul_mul_mux_113_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_96 <= MUX_s_1_2_2((MulIn_data_sva_133[96]), (mul_mul_mux_114_nl),
          and_dcpl_22);
      chn_mul_out_rsci_d_127 <= MUX_s_1_2_2((MulIn_data_sva_133[127]), (mul_mul_mux_115_nl),
          and_dcpl_22);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_out_rsci_d_22_1 <= 22'b0;
      chn_mul_out_rsci_d_30_23 <= 8'b0;
      chn_mul_out_rsci_d_54_33 <= 22'b0;
      chn_mul_out_rsci_d_62_55 <= 8'b0;
      chn_mul_out_rsci_d_86_65 <= 22'b0;
      chn_mul_out_rsci_d_94_87 <= 8'b0;
      chn_mul_out_rsci_d_118_97 <= 22'b0;
      chn_mul_out_rsci_d_126_119 <= 8'b0;
    end
    else if ( chn_mul_out_and_1_cse ) begin
      chn_mul_out_rsci_d_22_1 <= MUX1HOT_v_22_3_2((FpMul_8U_23U_o_mant_1_lpi_1_dfm_3[22:1]),
          (mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl),
          (MulIn_data_sva_133[22:1]), {(nor_3_nl) , asn_160 , asn_162});
      chn_mul_out_rsci_d_30_23 <= MUX1HOT_v_8_4_2((FpMul_8U_23U_FpMul_8U_23U_and_15_nl),
          FpMul_8U_23U_p_expo_1_sva_5, (MulIn_data_sva_133[30:23]), (mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl),
          {(and_358_nl) , (and_359_nl) , (or_839_nl) , asn_160});
      chn_mul_out_rsci_d_54_33 <= MUX1HOT_v_22_3_2((FpMul_8U_23U_o_mant_2_lpi_1_dfm_3[22:1]),
          (mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl),
          (MulIn_data_sva_133[54:33]), {(nor_2_nl) , asn_168 , asn_170});
      chn_mul_out_rsci_d_62_55 <= MUX1HOT_v_8_4_2((FpMul_8U_23U_FpMul_8U_23U_and_16_nl),
          FpMul_8U_23U_p_expo_2_sva_5, (MulIn_data_sva_133[62:55]), (mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl),
          {(and_356_nl) , (and_357_nl) , (or_838_nl) , asn_168});
      chn_mul_out_rsci_d_86_65 <= MUX1HOT_v_22_3_2((FpMul_8U_23U_o_mant_3_lpi_1_dfm_3[22:1]),
          (mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl),
          (MulIn_data_sva_133[86:65]), {(nor_1_nl) , asn_164 , asn_166});
      chn_mul_out_rsci_d_94_87 <= MUX1HOT_v_8_4_2((FpMul_8U_23U_FpMul_8U_23U_and_17_nl),
          FpMul_8U_23U_p_expo_3_sva_5, (MulIn_data_sva_133[94:87]), (mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl),
          {(and_354_nl) , (and_355_nl) , (or_837_nl) , asn_164});
      chn_mul_out_rsci_d_118_97 <= MUX1HOT_v_22_3_2((FpMul_8U_23U_o_mant_lpi_1_dfm_3[22:1]),
          (mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl),
          (MulIn_data_sva_133[118:97]), {(nor_6_nl) , asn_156 , asn_158});
      chn_mul_out_rsci_d_126_119 <= MUX1HOT_v_8_4_2((FpMul_8U_23U_FpMul_8U_23U_and_18_nl),
          FpMul_8U_23U_p_expo_sva_5, (MulIn_data_sva_133[126:119]), (mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl),
          {(and_352_nl) , (and_353_nl) , (or_836_nl) , asn_156});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_mul_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_24 | and_dcpl_26) ) begin
      reg_chn_mul_out_rsci_ld_core_psct_cse <= ~ and_dcpl_26;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_mul_op_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & (or_tmp_588 | chn_mul_op_rsci_ld_core_psct_mx0c1) ) begin
      chn_mul_op_rsci_ld_core_psct <= ~ chn_mul_op_rsci_ld_core_psct_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_591 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & not_tmp_2 ) begin
      IsZero_8U_23U_land_1_lpi_1_dfm_6 <= IsZero_8U_23U_land_1_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_132 <= 128'b0;
      io_read_cfg_mul_bypass_rsc_svs_st_4 <= 1'b0;
      mul_mul_land_1_lpi_1_dfm_5 <= 1'b0;
      mul_mul_land_2_lpi_1_dfm_5 <= 1'b0;
      mul_mul_land_3_lpi_1_dfm_5 <= 1'b0;
      mul_mul_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( MulIn_data_and_1_cse ) begin
      MulIn_data_sva_132 <= MulIn_data_sva_1;
      io_read_cfg_mul_bypass_rsc_svs_st_4 <= io_read_cfg_mul_bypass_rsc_svs_st_1;
      mul_mul_land_1_lpi_1_dfm_5 <= mul_mul_land_1_lpi_1_dfm_2;
      mul_mul_land_2_lpi_1_dfm_5 <= mul_mul_land_2_lpi_1_dfm_2;
      mul_mul_land_3_lpi_1_dfm_5 <= mul_mul_land_3_lpi_1_dfm_2;
      mul_mul_land_lpi_1_dfm_5 <= mul_mul_land_lpi_1_dfm_2;
      IsNaN_8U_23U_land_lpi_1_dfm_7 <= IsNaN_8U_23U_land_lpi_1_dfm_4;
      IsNaN_8U_23U_land_3_lpi_1_dfm_7 <= IsNaN_8U_23U_land_3_lpi_1_dfm_4;
      IsNaN_8U_23U_land_2_lpi_1_dfm_7 <= IsNaN_8U_23U_land_2_lpi_1_dfm_4;
      IsNaN_8U_23U_land_1_lpi_1_dfm_7 <= IsNaN_8U_23U_land_1_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & not_tmp_2
        ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp,
          IsZero_8U_23U_1_land_1_lpi_1_dfm_5, and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_0_lpi_1_dfm_2_30_0_1 <= 31'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( else_MulOp_data_and_8_cse ) begin
      else_MulOp_data_0_lpi_1_dfm_2_30_0_1 <= else_MulOp_data_0_lpi_1_dfm_mx1[30:0];
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= IsNaN_8U_23U_land_1_lpi_1_dfm_st_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & (~
        (mux_9_nl)) ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 <= 1'b0;
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0;
    end
    else if ( FpMul_8U_23U_oelse_1_and_4_cse ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 <= MUX_s_1_2_2(FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_6_lpi_1_dfm_st, and_dcpl_39);
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2 <= MUX_v_64_2_2(mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0,
          mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm, and_dcpl_38);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & not_tmp_8 ) begin
      IsZero_8U_23U_land_2_lpi_1_dfm_6 <= IsZero_8U_23U_land_2_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & not_tmp_8
        ) begin
      IsZero_8U_23U_1_land_2_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp,
          IsZero_8U_23U_1_land_2_lpi_1_dfm_5, and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_1_lpi_1_dfm_2_30_0_1 <= 31'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( else_MulOp_data_and_9_cse ) begin
      else_MulOp_data_1_lpi_1_dfm_2_30_0_1 <= else_MulOp_data_1_lpi_1_dfm_mx1[30:0];
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= IsNaN_8U_23U_land_2_lpi_1_dfm_st_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & (~
        (mux_14_nl)) ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 <= 1'b0;
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0;
    end
    else if ( FpMul_8U_23U_oelse_1_and_5_cse ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 <= MUX_s_1_2_2(FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_7_lpi_1_dfm_st, and_dcpl_39);
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2 <= MUX_v_64_2_2(mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0,
          mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm, and_dcpl_38);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & not_tmp_12 ) begin
      IsZero_8U_23U_land_3_lpi_1_dfm_6 <= IsZero_8U_23U_land_3_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & not_tmp_12
        ) begin
      IsZero_8U_23U_1_land_3_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp,
          IsZero_8U_23U_1_land_3_lpi_1_dfm_5, and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_2_lpi_1_dfm_2_30_0_1 <= 31'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( else_MulOp_data_and_10_cse ) begin
      else_MulOp_data_2_lpi_1_dfm_2_30_0_1 <= else_MulOp_data_2_lpi_1_dfm_mx1[30:0];
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= IsNaN_8U_23U_land_3_lpi_1_dfm_st_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & (~
        (mux_19_nl)) ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 <= 1'b0;
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0;
    end
    else if ( FpMul_8U_23U_oelse_1_and_6_cse ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 <= MUX_s_1_2_2(FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_8_lpi_1_dfm_st, and_dcpl_39);
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2 <= MUX_v_64_2_2(mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0,
          mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm, and_dcpl_38);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & not_tmp_15 ) begin
      IsZero_8U_23U_land_lpi_1_dfm_6 <= IsZero_8U_23U_land_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & not_tmp_15
        ) begin
      IsZero_8U_23U_1_land_lpi_1_dfm_6 <= MUX_s_1_2_2(IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp,
          IsZero_8U_23U_1_land_lpi_1_dfm_5, and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_3_lpi_1_dfm_2_30_0_1 <= 31'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( else_MulOp_data_and_11_cse ) begin
      else_MulOp_data_3_lpi_1_dfm_2_30_0_1 <= else_MulOp_data_3_lpi_1_dfm_mx1[30:0];
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= IsNaN_8U_23U_land_lpi_1_dfm_st_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse & (~
        (mux_24_nl)) ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
          <= MUX_s_1_2_2(mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= 1'b0;
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0;
    end
    else if ( FpMul_8U_23U_oelse_1_and_7_cse ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= MUX_s_1_2_2(FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0,
          FpMul_8U_23U_lor_1_lpi_1_dfm_st, and_dcpl_39);
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2 <= MUX_v_64_2_2(mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0,
          mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm, and_dcpl_38);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_land_lpi_1_dfm_st_4 <= 1'b0;
      mul_mul_land_3_lpi_1_dfm_st_4 <= 1'b0;
      mul_mul_land_2_lpi_1_dfm_st_4 <= 1'b0;
      mul_mul_land_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( mul_mul_aelse_and_cse ) begin
      mul_mul_land_lpi_1_dfm_st_4 <= mul_mul_land_lpi_1_dfm_st_1;
      mul_mul_land_3_lpi_1_dfm_st_4 <= mul_mul_land_3_lpi_1_dfm_st_1;
      mul_mul_land_2_lpi_1_dfm_st_4 <= mul_mul_land_2_lpi_1_dfm_st_1;
      mul_mul_land_1_lpi_1_dfm_st_4 <= mul_mul_land_1_lpi_1_dfm_st_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & ((or_74_cse & main_stage_v_2) | main_stage_v_3_mx0c1) )
        begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_133 <= 128'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
      mul_mul_land_lpi_1_dfm_6 <= 1'b0;
      mul_mul_land_3_lpi_1_dfm_6 <= 1'b0;
      mul_mul_land_2_lpi_1_dfm_6 <= 1'b0;
      mul_mul_land_1_lpi_1_dfm_6 <= 1'b0;
      io_read_cfg_mul_bypass_rsc_svs_5 <= 1'b0;
    end
    else if ( MulIn_data_and_2_cse ) begin
      MulIn_data_sva_133 <= MulIn_data_sva_132;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= IsNaN_8U_23U_land_1_lpi_1_dfm_7;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= IsNaN_8U_23U_land_2_lpi_1_dfm_7;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= IsNaN_8U_23U_land_3_lpi_1_dfm_7;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= IsNaN_8U_23U_land_lpi_1_dfm_7;
      mul_mul_land_lpi_1_dfm_6 <= mul_mul_land_lpi_1_dfm_5;
      mul_mul_land_3_lpi_1_dfm_6 <= mul_mul_land_3_lpi_1_dfm_5;
      mul_mul_land_2_lpi_1_dfm_6 <= mul_mul_land_2_lpi_1_dfm_5;
      mul_mul_land_1_lpi_1_dfm_6 <= mul_mul_land_1_lpi_1_dfm_5;
      io_read_cfg_mul_bypass_rsc_svs_5 <= io_read_cfg_mul_bypass_rsc_svs_st_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1 <= 32'b0;
      FpMul_8U_23U_mux_10_itm_4 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[31:0];
      FpMul_8U_23U_mux_10_itm_4 <= FpMul_8U_23U_mux_10_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1 <= 32'b0;
      FpMul_8U_23U_mux_23_itm_4 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[31:0];
      FpMul_8U_23U_mux_23_itm_4 <= FpMul_8U_23U_mux_23_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1 <= 32'b0;
      FpMul_8U_23U_mux_36_itm_4 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[31:0];
      FpMul_8U_23U_mux_36_itm_4 <= FpMul_8U_23U_mux_36_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1 <= 32'b0;
      FpMul_8U_23U_mux_49_itm_4 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse ) begin
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[31:0];
      FpMul_8U_23U_mux_49_itm_4 <= FpMul_8U_23U_mux_49_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_1_sva_5 <= 8'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse & (mux_42_nl)
        ) begin
      FpMul_8U_23U_p_expo_1_sva_5 <= MUX1HOT_v_8_4_2(FpMul_8U_23U_p_expo_1_sva_1_mx0w0,
          FpMul_8U_23U_p_expo_1_sva_1, (else_MulOp_data_0_lpi_1_dfm_2_30_0_1[30:23]),
          else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm, {and_dcpl_46 , and_dcpl_48
          , and_dcpl_50 , and_dcpl_51});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_44_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3
          <= MUX_s_1_2_2(mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1,
          FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2,
          and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_49_nl) ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_50_nl) ) begin
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= MUX_s_1_2_2((mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
          mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & (~ (mux_55_nl)) ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_cse ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[64];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2 <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_cse ) begin
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse & (mux_63_nl)
        ) begin
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2 <= MUX1HOT_v_23_4_2((else_MulOp_data_0_lpi_1_dfm_2_30_0_1[22:0]),
          else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm, (FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23]),
          mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1,
          {and_dcpl_50 , and_dcpl_51 , and_dcpl_46 , and_dcpl_48});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= 1'b0;
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_17_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & not_tmp_55 ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_7 <= FpMul_8U_23U_lor_6_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (~ mux_tmp_48) ) begin
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_1_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_66_nl) ) begin
      FpMantRNE_48U_24U_else_carry_1_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_1_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_1_sva, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse ) begin
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= MUX_s_1_2_2(mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0,
          mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm, and_dcpl_52);
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= MUX_s_1_2_2(mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0,
          mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm, and_dcpl_52);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_2_sva_5 <= 8'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse & (mux_74_nl)
        ) begin
      FpMul_8U_23U_p_expo_2_sva_5 <= MUX1HOT_v_8_4_2(FpMul_8U_23U_p_expo_2_sva_1_mx0w0,
          FpMul_8U_23U_p_expo_2_sva_1, (else_MulOp_data_1_lpi_1_dfm_2_30_0_1[30:23]),
          else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm, {and_dcpl_54 , and_dcpl_55
          , and_dcpl_57 , and_dcpl_58});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_76_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3
          <= MUX_s_1_2_2(mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1,
          FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2,
          and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_81_nl) ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_82_nl) ) begin
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= MUX_s_1_2_2((mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
          mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & (~ (mux_85_nl)) ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_1_cse ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[64];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2 <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_9_cse ) begin
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_12_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse & (mux_93_nl)
        ) begin
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2 <= MUX1HOT_v_23_4_2((else_MulOp_data_1_lpi_1_dfm_2_30_0_1[22:0]),
          else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm, (FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23]),
          mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1,
          {and_dcpl_57 , and_dcpl_58 , and_dcpl_54 , and_dcpl_55});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= 1'b0;
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_19_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & not_tmp_82 ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_7 <= FpMul_8U_23U_lor_7_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (~ mux_94_itm) ) begin
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_2_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_97_nl) ) begin
      FpMantRNE_48U_24U_else_carry_2_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_2_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_2_sva, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse ) begin
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= MUX_s_1_2_2(mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0,
          mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm, and_dcpl_52);
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= MUX_s_1_2_2(mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0,
          mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm, and_dcpl_52);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_3_sva_5 <= 8'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse & (mux_105_nl)
        ) begin
      FpMul_8U_23U_p_expo_3_sva_5 <= MUX1HOT_v_8_4_2(FpMul_8U_23U_p_expo_3_sva_1_mx0w0,
          FpMul_8U_23U_p_expo_3_sva_1, (else_MulOp_data_2_lpi_1_dfm_2_30_0_1[30:23]),
          else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm, {and_dcpl_60 , and_dcpl_61
          , and_dcpl_63 , and_dcpl_64});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_107_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3
          <= MUX_s_1_2_2(mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1,
          FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2,
          and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_112_nl) ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_113_nl) ) begin
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= MUX_s_1_2_2((mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
          mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & (~ (mux_116_nl)) ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_2_cse ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[64];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2 <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_11_cse ) begin
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_13_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse & (mux_124_nl)
        ) begin
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2 <= MUX1HOT_v_23_4_2((else_MulOp_data_2_lpi_1_dfm_2_30_0_1[22:0]),
          else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm, (FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23]),
          mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1,
          {and_dcpl_63 , and_dcpl_64 , and_dcpl_60 , and_dcpl_61});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= 1'b0;
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_21_cse ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & not_tmp_107 ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_7 <= FpMul_8U_23U_lor_8_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (~ mux_125_itm) ) begin
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_3_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_128_nl) ) begin
      FpMantRNE_48U_24U_else_carry_3_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_3_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_3_sva, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse ) begin
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= MUX_s_1_2_2(mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0,
          mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm, and_dcpl_52);
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= MUX_s_1_2_2(mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0,
          mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm, and_dcpl_52);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_sva_5 <= 8'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse & (mux_136_nl)
        ) begin
      FpMul_8U_23U_p_expo_sva_5 <= MUX1HOT_v_8_4_2(FpMul_8U_23U_p_expo_sva_1_mx0w0,
          FpMul_8U_23U_p_expo_sva_1, (else_MulOp_data_3_lpi_1_dfm_2_30_0_1[30:23]),
          else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm, {and_dcpl_66 , and_dcpl_67
          , and_dcpl_69 , and_dcpl_70});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_138_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3
          <= MUX_s_1_2_2(mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1,
          FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2,
          and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_143_nl) ) begin
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0,
          FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (~ (mux_147_nl)) ) begin
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= MUX_s_1_2_2((mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]),
          mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & (~ (mux_149_nl)) ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
          <= mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_3_cse ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_lpi_1_dfm_6;
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1 <= IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[64];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2 <= 1'b0;
    end
    else if ( FpMantRNE_48U_24U_else_and_13_cse ) begin
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2 <= MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0,
          FpMul_8U_23U_FpMul_8U_23U_and_14_itm, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse & (mux_156_nl)
        ) begin
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2 <= MUX1HOT_v_23_4_2((else_MulOp_data_3_lpi_1_dfm_2_30_0_1[22:0]),
          else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm, (FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23]),
          mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1,
          {and_dcpl_69 , and_dcpl_70 , and_dcpl_66 , and_dcpl_67});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= 1'b0;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_23_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_lpi_1_dfm_st_4;
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_23) & not_tmp_130 ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_7 <= FpMul_8U_23U_lor_1_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (~ mux_tmp_140) ) begin
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2 <= FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_48U_24U_else_carry_sva_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse
        & (mux_159_nl) ) begin
      FpMantRNE_48U_24U_else_carry_sva_2 <= MUX_s_1_2_2(FpMantRNE_48U_24U_else_carry_sva_mx0w0,
          FpMantRNE_48U_24U_else_carry_sva, and_dcpl_47);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse ) begin
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= MUX_s_1_2_2(mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0,
          mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm, and_dcpl_52);
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= MUX_s_1_2_2(mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0,
          mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm, and_dcpl_52);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_land_lpi_1_dfm_st_5 <= 1'b0;
      mul_mul_land_3_lpi_1_dfm_st_5 <= 1'b0;
      mul_mul_land_2_lpi_1_dfm_st_5 <= 1'b0;
      mul_mul_land_1_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( mul_mul_aelse_and_12_cse ) begin
      mul_mul_land_lpi_1_dfm_st_5 <= mul_mul_land_lpi_1_dfm_st_4;
      mul_mul_land_3_lpi_1_dfm_st_5 <= mul_mul_land_3_lpi_1_dfm_st_4;
      mul_mul_land_2_lpi_1_dfm_st_5 <= mul_mul_land_2_lpi_1_dfm_st_4;
      mul_mul_land_1_lpi_1_dfm_st_5 <= mul_mul_land_1_lpi_1_dfm_st_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_587 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      MulIn_data_sva_1 <= 128'b0;
      io_read_cfg_mul_bypass_rsc_svs_st_1 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
      mul_mul_land_1_lpi_1_dfm_2 <= 1'b0;
      mul_mul_land_2_lpi_1_dfm_2 <= 1'b0;
      mul_mul_land_3_lpi_1_dfm_2 <= 1'b0;
      mul_mul_land_lpi_1_dfm_2 <= 1'b0;
      cfg_truncate_1_sva_1 <= 10'b0;
    end
    else if ( MulIn_data_and_cse ) begin
      MulIn_data_sva_1 <= chn_mul_in_rsci_d_mxwt;
      io_read_cfg_mul_bypass_rsc_svs_st_1 <= cfg_mul_bypass_rsci_d;
      IsNaN_8U_23U_land_1_lpi_1_dfm_4 <= IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
      mul_mul_land_1_lpi_1_dfm_2 <= mul_mul_land_1_lpi_1_dfm_mx1w0;
      mul_mul_land_2_lpi_1_dfm_2 <= mul_mul_land_2_lpi_1_dfm_mx1w0;
      mul_mul_land_3_lpi_1_dfm_2 <= mul_mul_land_3_lpi_1_dfm_mx1w0;
      mul_mul_land_lpi_1_dfm_2 <= mul_mul_land_lpi_1_dfm_mx1w0;
      cfg_truncate_1_sva_1 <= cfg_truncate_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_1 <= 1'b0;
      IsZero_8U_23U_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_24_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_1_lpi_1_dfm_st, and_dcpl_6);
      IsZero_8U_23U_land_1_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0,
          IsZero_8U_23U_land_1_lpi_1_dfm, and_dcpl_6);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_op_1_sva_1 <= 32'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_cse & and_20_tmp & (~(or_tmp_461 | cfg_mul_src_rsci_d))
        ) begin
      cfg_mul_op_1_sva_1 <= cfg_mul_op_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_1_sva_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_cse & and_20_tmp & (~ or_tmp_461) ) begin
      cfg_mul_src_1_sva_1 <= cfg_mul_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_1 <= 1'b0;
      IsZero_8U_23U_land_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_25_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_2_lpi_1_dfm_st, and_dcpl_6);
      IsZero_8U_23U_land_2_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0,
          IsZero_8U_23U_land_2_lpi_1_dfm, and_dcpl_6);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_1 <= 1'b0;
      IsZero_8U_23U_land_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_26_cse ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_3_lpi_1_dfm_st, and_dcpl_6);
      IsZero_8U_23U_land_3_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0,
          IsZero_8U_23U_land_3_lpi_1_dfm, and_dcpl_6);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_1 <= 1'b0;
      IsZero_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_27_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_1 <= MUX_s_1_2_2(IsNaN_8U_23U_land_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_land_lpi_1_dfm_st, and_dcpl_6);
      IsZero_8U_23U_land_lpi_1_dfm_4 <= MUX_s_1_2_2(IsZero_8U_23U_land_lpi_1_dfm_mx1w0,
          IsZero_8U_23U_land_lpi_1_dfm, and_dcpl_6);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_land_lpi_1_dfm_st_1 <= 1'b0;
      mul_mul_land_3_lpi_1_dfm_st_1 <= 1'b0;
      mul_mul_land_2_lpi_1_dfm_st_1 <= 1'b0;
      mul_mul_land_1_lpi_1_dfm_st_1 <= 1'b0;
    end
    else if ( mul_mul_aelse_and_19_cse ) begin
      mul_mul_land_lpi_1_dfm_st_1 <= mul_mul_land_lpi_1_dfm_mx1w0;
      mul_mul_land_3_lpi_1_dfm_st_1 <= mul_mul_land_3_lpi_1_dfm_mx1w0;
      mul_mul_land_2_lpi_1_dfm_st_1 <= mul_mul_land_2_lpi_1_dfm_mx1w0;
      mul_mul_land_1_lpi_1_dfm_st_1 <= mul_mul_land_1_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_1_sva_st_1 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_27 & (fsm_output[1])) | cfg_mul_src_1_sva_st_1_mx0c1)
        ) begin
      cfg_mul_src_1_sva_st_1 <= MUX_s_1_2_2(cfg_mul_src_rsci_d, cfg_mul_src_1_sva_st,
          cfg_mul_src_1_sva_st_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_22) & (mux_185_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2
          <= mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_27) & (mux_187_nl) ) begin
      mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_1_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm <= 1'b0;
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_cse ) begin
      FpMul_8U_23U_p_expo_1_sva_1 <= FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0;
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm <= 8'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | or_dcpl_23 | (~ (cfg_precision[1])) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_4))
        ) begin
      else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm <= else_MulOp_data_0_lpi_1_dfm_2_30_0_1[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm <= 23'b0;
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
      FpMantRNE_48U_24U_else_carry_1_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_itm <= 1'b0;
    end
    else if ( else_MulOp_data_and_1_cse ) begin
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm <= else_MulOp_data_0_lpi_1_dfm_2_30_0_1[22:0];
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st <= mul_mul_1_FpMantRNE_48U_24U_else_and_tmp;
      FpMantRNE_48U_24U_else_carry_1_sva <= FpMantRNE_48U_24U_else_carry_1_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_itm <= FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_cse ) begin
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_37) & (mux_189_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2
          <= mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_40) & (mux_191_nl) ) begin
      mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_2_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm <= 1'b0;
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_1_cse ) begin
      FpMul_8U_23U_p_expo_2_sva_1 <= FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0;
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm <= 8'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | mul_mul_land_2_lpi_1_dfm_st_4 | IsNaN_8U_23U_land_2_lpi_1_dfm_st_4
        | or_27_cse)) ) begin
      else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm <= else_MulOp_data_1_lpi_1_dfm_2_30_0_1[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm <= 23'b0;
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
      FpMantRNE_48U_24U_else_carry_2_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm <= 1'b0;
    end
    else if ( else_MulOp_data_and_3_cse ) begin
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm <= else_MulOp_data_1_lpi_1_dfm_2_30_0_1[22:0];
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st <= mul_mul_2_FpMantRNE_48U_24U_else_and_tmp;
      FpMantRNE_48U_24U_else_carry_2_sva <= FpMantRNE_48U_24U_else_carry_2_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm <= FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse ) begin
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_50) & (mux_193_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2
          <= mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_53) & (mux_195_nl) ) begin
      mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_3_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm <= 1'b0;
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_2_cse ) begin
      FpMul_8U_23U_p_expo_3_sva_1 <= FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0;
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm <= 8'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | mul_mul_land_3_lpi_1_dfm_st_4 | IsNaN_8U_23U_land_3_lpi_1_dfm_st_4
        | or_27_cse)) ) begin
      else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm <= else_MulOp_data_2_lpi_1_dfm_2_30_0_1[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm <= 23'b0;
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
      FpMantRNE_48U_24U_else_carry_3_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm <= 1'b0;
    end
    else if ( else_MulOp_data_and_5_cse ) begin
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm <= else_MulOp_data_2_lpi_1_dfm_2_30_0_1[22:0];
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st <= mul_mul_3_FpMantRNE_48U_24U_else_and_tmp;
      FpMantRNE_48U_24U_else_carry_3_sva <= FpMantRNE_48U_24U_else_carry_3_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm <= FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse ) begin
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_63) & (mux_197_nl) ) begin
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2
          <= mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= 23'b0;
    end
    else if ( core_wen & (~ or_dcpl_66) & (mux_201_nl) ) begin
      mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1
          <= FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_expo_sva_1 <= 8'b0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm <= 1'b0;
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    end
    else if ( FpMul_8U_23U_p_expo_and_3_cse ) begin
      FpMul_8U_23U_p_expo_sva_1 <= FpMul_8U_23U_p_expo_sva_1_mx0w0;
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm <= FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0;
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm <= 8'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | mul_mul_land_lpi_1_dfm_st_4 | IsNaN_8U_23U_land_lpi_1_dfm_st_4
        | or_27_cse)) ) begin
      else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm <= else_MulOp_data_3_lpi_1_dfm_2_30_0_1[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm <= 23'b0;
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
      FpMantRNE_48U_24U_else_carry_sva <= 1'b0;
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm <= 1'b0;
    end
    else if ( else_MulOp_data_and_7_cse ) begin
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm <= else_MulOp_data_3_lpi_1_dfm_2_30_0_1[22:0];
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st <= mul_mul_4_FpMantRNE_48U_24U_else_and_tmp;
      FpMantRNE_48U_24U_else_carry_sva <= FpMantRNE_48U_24U_else_carry_sva_mx0w0;
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm <= FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    end
    else if ( IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse ) begin
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (mux_203_nl) ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_6 <= (FpMul_8U_23U_oelse_1_mux_20_nl) & (~ and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & (~(mul_mul_land_1_lpi_1_dfm_2 | mul_mul_land_1_lpi_1_dfm_st_1
        | io_read_cfg_mul_bypass_rsc_svs_st_1)) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_10_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_135_rgt | mul_mul_if_and_6_rgt | mul_mul_if_and_7_rgt)
        & (mux_207_nl) ) begin
      FpMul_8U_23U_mux_10_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_1[31]), (mul_mul_1_FpMul_8U_23U_xor_nl),
          (else_MulOp_data_0_lpi_1_dfm_mx1[31]), {and_135_rgt , mul_mul_if_and_6_rgt
          , mul_mul_if_and_7_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (mux_209_nl) ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_6 <= (FpMul_8U_23U_oelse_1_mux_21_nl) & (~ and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & (~(mul_mul_land_2_lpi_1_dfm_2 | mul_mul_land_2_lpi_1_dfm_st_1
        | io_read_cfg_mul_bypass_rsc_svs_st_1)) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_23_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_137_rgt | mul_mul_if_and_4_rgt | mul_mul_if_and_5_rgt)
        & (mux_213_nl) ) begin
      FpMul_8U_23U_mux_23_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_1[63]), (mul_mul_2_FpMul_8U_23U_xor_nl),
          (else_MulOp_data_1_lpi_1_dfm_mx1[31]), {and_137_rgt , mul_mul_if_and_4_rgt
          , mul_mul_if_and_5_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (mux_215_nl) ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_6 <= (FpMul_8U_23U_oelse_1_mux_22_nl) & (~ and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & (~(mul_mul_land_3_lpi_1_dfm_2 | mul_mul_land_3_lpi_1_dfm_st_1
        | io_read_cfg_mul_bypass_rsc_svs_st_1)) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_36_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_139_rgt | mul_mul_if_and_2_rgt | mul_mul_if_and_3_rgt)
        & (mux_219_nl) ) begin
      FpMul_8U_23U_mux_36_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_1[95]), (mul_mul_3_FpMul_8U_23U_xor_nl),
          (else_MulOp_data_2_lpi_1_dfm_mx1[31]), {and_139_rgt , mul_mul_if_and_2_rgt
          , mul_mul_if_and_3_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (mux_221_nl) ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_6 <= (FpMul_8U_23U_oelse_1_mux_23_nl) & (~ and_dcpl_39);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & and_18_tmp & (~(mul_mul_land_lpi_1_dfm_2 | mul_mul_land_lpi_1_dfm_st_1
        | io_read_cfg_mul_bypass_rsc_svs_st_1)) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_mux_49_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_141_rgt | mul_mul_if_and_rgt | mul_mul_if_and_1_rgt)
        & (mux_225_nl) ) begin
      FpMul_8U_23U_mux_49_itm_3 <= MUX1HOT_s_1_3_2((MulIn_data_sva_1[127]), (mul_mul_4_FpMul_8U_23U_xor_nl),
          (else_MulOp_data_3_lpi_1_dfm_mx1[31]), {and_141_rgt , mul_mul_if_and_rgt
          , mul_mul_if_and_1_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_1_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | mul_mul_land_1_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3
        | or_27_cse)) & mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_1_sva <= mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          1'b0;
    end
    else if ( core_wen & ((nor_118_cse & and_dcpl_38) | and_146_rgt) & (~ mux_7_itm)
        ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          MUX_s_1_2_2(mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_146_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_truncate_1_sva_3 <= 10'b0;
    end
    else if ( core_wen & and_18_tmp & (~((mul_mul_land_2_lpi_1_dfm_st_1 & mul_mul_land_lpi_1_dfm_st_1
        & mul_mul_land_1_lpi_1_dfm_st_1 & mul_mul_land_3_lpi_1_dfm_st_1) | io_read_cfg_mul_bypass_rsc_svs_st_1))
        ) begin
      cfg_truncate_1_sva_3 <= cfg_truncate_1_sva_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_2_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | or_tmp_252 | or_27_cse)) & mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_2_sva <= mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          1'b0;
    end
    else if ( core_wen & ((nor_117_cse & and_dcpl_38) | and_150_rgt) & (~ mux_12_itm)
        ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          MUX_s_1_2_2(mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_150_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_3_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | or_tmp_332 | or_27_cse)) & mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_3_sva <= mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          1'b0;
    end
    else if ( core_wen & ((nor_116_cse & and_dcpl_38) | and_154_rgt) & (~ mux_17_itm)
        ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          MUX_s_1_2_2(mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_154_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_p_mant_p1_sva <= 48'b0;
    end
    else if ( core_wen & (~(or_dcpl_26 | mul_mul_land_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
        | or_27_cse)) & mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3
        ) begin
      FpMul_8U_23U_p_mant_p1_sva <= mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          1'b0;
    end
    else if ( core_wen & ((nor_115_cse & and_dcpl_38) | and_158_rgt) & (~ mux_22_itm)
        ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <=
          MUX_s_1_2_2(mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1, mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs,
          and_158_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_99) & (~ (mux_164_nl)) ) begin
      IsZero_8U_23U_1_land_1_lpi_1_dfm_5 <= IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_99 | (fsm_output[0]))) ) begin
      FpMul_8U_23U_lor_6_lpi_1_dfm_st <= FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_102) & (~ (mux_172_nl)) ) begin
      IsZero_8U_23U_1_land_2_lpi_1_dfm_5 <= IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_102 | (fsm_output[0]))) ) begin
      FpMul_8U_23U_lor_7_lpi_1_dfm_st <= FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_105) & (~ (mux_177_nl)) ) begin
      IsZero_8U_23U_1_land_3_lpi_1_dfm_5 <= IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_105 | (fsm_output[0]))) ) begin
      FpMul_8U_23U_lor_8_lpi_1_dfm_st <= FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_8U_23U_1_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_108) & (~ (mux_182_nl)) ) begin
      IsZero_8U_23U_1_land_lpi_1_dfm_5 <= IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_108 | (fsm_output[0]))) ) begin
      FpMul_8U_23U_lor_1_lpi_1_dfm_st <= FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_4_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st <= IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_land_1_lpi_1_dfm <= IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_5_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_st <= IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_land_2_lpi_1_dfm <= IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_6_cse ) begin
      IsNaN_8U_23U_land_3_lpi_1_dfm_st <= IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_land_3_lpi_1_dfm <= IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st <= 1'b0;
      IsZero_8U_23U_land_lpi_1_dfm <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_7_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st <= IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
      IsZero_8U_23U_land_lpi_1_dfm <= IsZero_8U_23U_land_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_mul_src_1_sva_st <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_8 | (fsm_output[0]))) ) begin
      cfg_mul_src_1_sva_st <= cfg_mul_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_75 | IsZero_8U_23U_land_1_lpi_1_dfm_4 | io_read_cfg_mul_bypass_rsc_svs_st_1
        | mul_mul_land_1_lpi_1_dfm_st_1 | (cfg_precision[0]) | or_dcpl_96 | (fsm_output[0])))
        ) begin
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0;
    end
    else if ( core_wen & (~(or_dcpl_125 | mul_mul_land_1_lpi_1_dfm_st_1 | (~ and_18_tmp)
        | (fsm_output[0]))) ) begin
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm <= mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_81 | IsZero_8U_23U_land_2_lpi_1_dfm_4 | io_read_cfg_mul_bypass_rsc_svs_st_1
        | mul_mul_land_2_lpi_1_dfm_st_1 | (cfg_precision[0]) | or_dcpl_96 | (fsm_output[0])))
        ) begin
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0;
    end
    else if ( core_wen & (~(or_dcpl_125 | mul_mul_land_2_lpi_1_dfm_st_1 | (~ and_18_tmp)
        | (fsm_output[0]))) ) begin
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm <= mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_87 | IsZero_8U_23U_land_3_lpi_1_dfm_4 | io_read_cfg_mul_bypass_rsc_svs_st_1
        | mul_mul_land_3_lpi_1_dfm_st_1 | (cfg_precision[0]) | or_dcpl_96 | (fsm_output[0])))
        ) begin
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0;
    end
    else if ( core_wen & (~(or_dcpl_125 | mul_mul_land_3_lpi_1_dfm_st_1 | (~ and_18_tmp)
        | (fsm_output[0]))) ) begin
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm <= mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_93 | mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1
        | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_lpi_1_dfm_st_1 | (cfg_precision[0])
        | or_dcpl_96 | (fsm_output[0]))) ) begin
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0;
    end
    else if ( core_wen & (~(or_dcpl_125 | mul_mul_land_lpi_1_dfm_st_1 | (~ and_18_tmp)
        | (fsm_output[0]))) ) begin
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm <= mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
    end
  end
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[0]) |
      IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva)) | IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva);
  assign mul_mul_else_mux_26_nl = MUX_s_1_2_2((FpMul_8U_23U_o_mant_1_lpi_1_dfm_3[0]),
      (mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_108_nl = MUX_s_1_2_2((mul_mul_else_mux_26_nl), (MulIn_data_sva_133[0]),
      mul_mul_land_1_lpi_1_dfm_6);
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[31]) |
      IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva)) | IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva);
  assign mul_mul_else_mux_23_nl = MUX_s_1_2_2(FpMul_8U_23U_mux_10_itm_4, (mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_109_nl = MUX_s_1_2_2((mul_mul_else_mux_23_nl), (MulIn_data_sva_133[31]),
      mul_mul_land_1_lpi_1_dfm_6);
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[0]) |
      IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva)) | IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva);
  assign mul_mul_else_mux_53_nl = MUX_s_1_2_2((FpMul_8U_23U_o_mant_2_lpi_1_dfm_3[0]),
      (mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_110_nl = MUX_s_1_2_2((mul_mul_else_mux_53_nl), (MulIn_data_sva_133[32]),
      mul_mul_land_2_lpi_1_dfm_6);
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[31]) |
      IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva)) | IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva);
  assign mul_mul_else_mux_50_nl = MUX_s_1_2_2(FpMul_8U_23U_mux_23_itm_4, (mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_111_nl = MUX_s_1_2_2((mul_mul_else_mux_50_nl), (MulIn_data_sva_133[63]),
      mul_mul_land_2_lpi_1_dfm_6);
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[0]) |
      IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva)) | IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva);
  assign mul_mul_else_mux_80_nl = MUX_s_1_2_2((FpMul_8U_23U_o_mant_3_lpi_1_dfm_3[0]),
      (mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_112_nl = MUX_s_1_2_2((mul_mul_else_mux_80_nl), (MulIn_data_sva_133[64]),
      mul_mul_land_3_lpi_1_dfm_6);
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[31]) |
      IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva)) | IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva);
  assign mul_mul_else_mux_77_nl = MUX_s_1_2_2(FpMul_8U_23U_mux_36_itm_4, (mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_113_nl = MUX_s_1_2_2((mul_mul_else_mux_77_nl), (MulIn_data_sva_133[95]),
      mul_mul_land_3_lpi_1_dfm_6);
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[0]) | IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva))
      | IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva);
  assign mul_mul_else_mux_107_nl = MUX_s_1_2_2((FpMul_8U_23U_o_mant_lpi_1_dfm_3[0]),
      (mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_114_nl = MUX_s_1_2_2((mul_mul_else_mux_107_nl), (MulIn_data_sva_133[96]),
      mul_mul_land_lpi_1_dfm_6);
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl
      = ~((~((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[31]) | IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva))
      | IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva);
  assign mul_mul_else_mux_104_nl = MUX_s_1_2_2(FpMul_8U_23U_mux_49_itm_4, (mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      mul_mul_else_unequal_tmp_1);
  assign mul_mul_mux_115_nl = MUX_s_1_2_2((mul_mul_else_mux_104_nl), (MulIn_data_sva_133[127]),
      mul_mul_land_lpi_1_dfm_6);
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~(MUX_v_22_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[22:1]),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva));
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl
      = ~(MUX_v_22_2_2((mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva));
  assign nor_3_nl = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_1_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5);
  assign FpMul_8U_23U_oelse_2_not_4_nl = ~ FpMul_8U_23U_lor_9_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_15_nl = MUX_v_8_2_2(8'b00000000, FpMul_8U_23U_o_expo_1_lpi_1_dfm,
      (FpMul_8U_23U_oelse_2_not_4_nl));
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~(MUX_v_8_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[30:23]),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva));
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl
      = ~(MUX_v_8_2_2((mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva));
  assign and_358_nl = (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7) & mul_mul_and_m1c;
  assign and_359_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & mul_mul_and_m1c;
  assign or_839_nl = (IsNaN_8U_23U_land_1_lpi_1_dfm_8 & mul_mul_mul_mul_nor_m1c &
      (~ io_read_cfg_mul_bypass_rsc_svs_5)) | asn_162;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~(MUX_v_22_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[22:1]),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva));
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl
      = ~(MUX_v_22_2_2((mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva));
  assign nor_2_nl = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_2_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5);
  assign FpMul_8U_23U_oelse_2_not_5_nl = ~ FpMul_8U_23U_lor_10_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_16_nl = MUX_v_8_2_2(8'b00000000, FpMul_8U_23U_o_expo_2_lpi_1_dfm,
      (FpMul_8U_23U_oelse_2_not_5_nl));
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~(MUX_v_8_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[30:23]),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva));
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl
      = ~(MUX_v_8_2_2((mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva));
  assign and_356_nl = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) & mul_mul_and_17_m1c;
  assign and_357_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & mul_mul_and_17_m1c;
  assign or_838_nl = (IsNaN_8U_23U_land_2_lpi_1_dfm_8 & mul_mul_mul_mul_nor_2_m1c
      & (~ io_read_cfg_mul_bypass_rsc_svs_5)) | asn_170;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~(MUX_v_22_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[22:1]),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva));
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl
      = ~(MUX_v_22_2_2((mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva));
  assign nor_1_nl = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_3_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5);
  assign FpMul_8U_23U_oelse_2_not_6_nl = ~ FpMul_8U_23U_lor_11_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_17_nl = MUX_v_8_2_2(8'b00000000, FpMul_8U_23U_o_expo_3_lpi_1_dfm,
      (FpMul_8U_23U_oelse_2_not_6_nl));
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~(MUX_v_8_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[30:23]),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva));
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl
      = ~(MUX_v_8_2_2((mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva));
  assign and_354_nl = (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7) & mul_mul_and_19_m1c;
  assign and_355_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & mul_mul_and_19_m1c;
  assign or_837_nl = (IsNaN_8U_23U_land_3_lpi_1_dfm_8 & mul_mul_mul_mul_nor_4_m1c
      & (~ io_read_cfg_mul_bypass_rsc_svs_5)) | asn_166;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~(MUX_v_22_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[22:1]),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva));
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl
      = ~(MUX_v_22_2_2((mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl),
      22'b1111111111111111111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva));
  assign nor_6_nl = ~(mul_mul_else_unequal_tmp_1 | mul_mul_land_lpi_1_dfm_6 | io_read_cfg_mul_bypass_rsc_svs_5);
  assign FpMul_8U_23U_oelse_2_not_7_nl = ~ FpMul_8U_23U_lor_2_lpi_1_dfm;
  assign FpMul_8U_23U_FpMul_8U_23U_and_18_nl = MUX_v_8_2_2(8'b00000000, FpMul_8U_23U_o_expo_lpi_1_dfm,
      (FpMul_8U_23U_oelse_2_not_7_nl));
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~(MUX_v_8_2_2((IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[30:23]),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva));
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl
      = ~(MUX_v_8_2_2((mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl),
      8'b11111111, IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva));
  assign and_352_nl = (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7) & mul_mul_and_21_m1c;
  assign and_353_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & mul_mul_and_21_m1c;
  assign or_836_nl = (IsNaN_8U_23U_land_lpi_1_dfm_8 & mul_mul_mul_mul_nor_6_m1c &
      (~ io_read_cfg_mul_bypass_rsc_svs_5)) | asn_158;
  assign or_28_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st | mul_mul_land_1_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign mux_8_nl = MUX_s_1_2_2(or_tmp_12, (or_28_nl), or_27_cse);
  assign or_31_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | mul_mul_land_1_lpi_1_dfm_st_4
      | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2);
  assign mux_9_nl = MUX_s_1_2_2((or_31_nl), (mux_8_nl), and_18_tmp);
  assign or_42_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st | mul_mul_land_2_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign mux_13_nl = MUX_s_1_2_2(or_tmp_26, (or_42_nl), or_27_cse);
  assign or_45_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | mul_mul_land_2_lpi_1_dfm_st_4
      | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2);
  assign mux_14_nl = MUX_s_1_2_2((or_45_nl), (mux_13_nl), and_18_tmp);
  assign or_56_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st | mul_mul_land_3_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_40, (or_56_nl), or_27_cse);
  assign or_59_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | mul_mul_land_3_lpi_1_dfm_st_4
      | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2);
  assign mux_19_nl = MUX_s_1_2_2((or_59_nl), (mux_18_nl), and_18_tmp);
  assign or_67_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st | mul_mul_land_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign mux_23_nl = MUX_s_1_2_2(or_tmp_51, (or_67_nl), or_27_cse);
  assign or_70_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ reg_chn_mul_out_rsci_ld_core_psct_cse)
      | chn_mul_out_rsci_bawt | mul_mul_land_lpi_1_dfm_st_4 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | (~ main_stage_v_2);
  assign mux_24_nl = MUX_s_1_2_2((or_70_nl), (mux_23_nl), and_18_tmp);
  assign nor_299_nl = ~(IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5);
  assign or_142_nl = nor_301_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5;
  assign or_143_nl = (~ FpMul_8U_23U_lor_6_lpi_1_dfm_6) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5;
  assign mux_35_nl = MUX_s_1_2_2((or_143_nl), (or_142_nl), mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_36_nl = MUX_s_1_2_2((mux_35_nl), or_tmp_123, mul_mul_1_FpMantRNE_48U_24U_else_and_tmp);
  assign or_147_nl = (~ or_tmp_128) | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5;
  assign mux_37_nl = MUX_s_1_2_2((or_147_nl), or_tmp_123, mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st);
  assign or_831_nl = (~((FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2
      & mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm) | FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm))
      | (mux_37_nl);
  assign mux_38_nl = MUX_s_1_2_2((or_831_nl), (mux_36_nl), nor_20_cse);
  assign nor_300_nl = ~(FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (mux_38_nl));
  assign mux_39_nl = MUX_s_1_2_2((nor_300_nl), (nor_299_nl), IsNaN_8U_23U_1_land_1_lpi_1_dfm_6);
  assign and_344_nl = (~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | (~ main_stage_v_2))) & (mux_39_nl);
  assign nor_304_nl = ~((~ or_tmp_133) | mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2
      | (~ or_tmp_132));
  assign mux_40_nl = MUX_s_1_2_2((nor_304_nl), or_tmp_132, mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2);
  assign or_153_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | (~(mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & (mux_40_nl)));
  assign mux_41_nl = MUX_s_1_2_2((or_153_nl), IsNaN_8U_23U_land_1_lpi_1_dfm_st_5,
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7);
  assign nor_303_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_8 | mul_mul_land_1_lpi_1_dfm_st_5 | (mux_41_nl));
  assign mux_42_nl = MUX_s_1_2_2((nor_303_nl), (and_344_nl), or_74_cse);
  assign nor_296_nl = ~((~ (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_1_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | nand_48_cse);
  assign nor_297_nl = ~((~ mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3
      | nand_48_cse);
  assign mux_43_nl = MUX_s_1_2_2((nor_297_nl), (nor_296_nl), nor_20_cse);
  assign nor_298_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | (~(mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2)));
  assign mux_44_nl = MUX_s_1_2_2((nor_298_nl), (mux_43_nl), or_74_cse);
  assign or_165_nl = nor_301_cse | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5;
  assign or_166_nl = (~ FpMul_8U_23U_lor_6_lpi_1_dfm_6) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5;
  assign mux_45_nl = MUX_s_1_2_2((or_166_nl), (or_165_nl), mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_46_nl = MUX_s_1_2_2((mux_45_nl), or_tmp_146, mul_mul_1_FpMantRNE_48U_24U_else_and_tmp);
  assign or_169_nl = (~ or_tmp_128) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5;
  assign mux_47_nl = MUX_s_1_2_2((or_169_nl), or_tmp_146, mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st);
  assign mux_48_nl = MUX_s_1_2_2((mux_47_nl), (mux_46_nl), nor_20_cse);
  assign nor_292_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (mux_48_nl));
  assign nor_294_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_8 | mul_mul_land_1_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_7
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | (~(mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & (mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 | (~((~ or_tmp_133) | mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2))))));
  assign mux_49_nl = MUX_s_1_2_2((nor_294_nl), (nor_292_nl), or_74_cse);
  assign nor_290_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | nand_48_cse);
  assign nor_291_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign mux_50_nl = MUX_s_1_2_2((nor_291_nl), (nor_290_nl), or_74_cse);
  assign or_181_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | mul_mul_land_1_lpi_1_dfm_st_5
      | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt | io_read_cfg_mul_bypass_rsc_svs_5
      | (~ main_stage_v_3);
  assign or_185_nl = mul_mul_land_1_lpi_1_dfm_st_4 | or_tmp_167;
  assign mux_54_nl = MUX_s_1_2_2(mux_tmp_48, (or_185_nl), FpMul_8U_23U_lor_6_lpi_1_dfm_st_4);
  assign mux_55_nl = MUX_s_1_2_2((mux_54_nl), (or_181_nl), FpMul_8U_23U_lor_6_lpi_1_dfm_st_3);
  assign nor_276_nl = ~(nor_277_cse | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5);
  assign nor_278_nl = ~((FpMul_8U_23U_p_mant_p1_1_sva[47]) | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5);
  assign mux_60_nl = MUX_s_1_2_2((nor_278_nl), (nor_276_nl), nor_31_cse);
  assign nand_15_nl = ~(mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_60_nl));
  assign or_210_nl = (~ FpMul_8U_23U_FpMul_8U_23U_and_itm) | IsNaN_8U_23U_land_1_lpi_1_dfm_7
      | mul_mul_land_1_lpi_1_dfm_5;
  assign mux_61_nl = MUX_s_1_2_2((or_210_nl), (nand_15_nl), nor_20_cse);
  assign or_211_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_6 | (mux_61_nl);
  assign mux_62_nl = MUX_s_1_2_2((or_211_nl), or_tmp_123, IsNaN_8U_23U_1_land_1_lpi_1_dfm_6);
  assign nor_275_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (mux_62_nl));
  assign nor_279_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_8 | mul_mul_land_1_lpi_1_dfm_st_5 | (~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_7
      | (~(nor_282_cse | FpMul_8U_23U_lor_6_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_itm_2))))));
  assign mux_63_nl = MUX_s_1_2_2((nor_279_nl), (nor_275_nl), or_74_cse);
  assign nor_269_nl = ~(nor_277_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | FpMul_8U_23U_lor_6_lpi_1_dfm_6 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6
      | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5);
  assign nor_271_nl = ~((FpMul_8U_23U_p_mant_p1_1_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_1_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_6_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5);
  assign mux_64_nl = MUX_s_1_2_2((nor_271_nl), (nor_269_nl), nor_31_cse);
  assign and_343_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_64_nl);
  assign nor_272_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_1_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_6_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5);
  assign mux_65_nl = MUX_s_1_2_2((nor_272_nl), (and_343_nl), nor_20_cse);
  assign nor_273_nl = ~(nor_282_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5
      | mul_mul_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_8 | mul_mul_land_1_lpi_1_dfm_st_5
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 | FpMul_8U_23U_lor_6_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_itm_2));
  assign mux_66_nl = MUX_s_1_2_2((nor_273_nl), (mux_65_nl), or_74_cse);
  assign or_227_nl = IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 | IsNaN_8U_23U_land_2_lpi_1_dfm_7
      | mul_mul_land_2_lpi_1_dfm_5;
  assign or_230_nl = nor_264_cse | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign or_231_nl = (~ FpMul_8U_23U_lor_7_lpi_1_dfm_6) | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3
      | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign mux_67_nl = MUX_s_1_2_2((or_231_nl), (or_230_nl), mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_68_nl = MUX_s_1_2_2((mux_67_nl), or_tmp_211, mul_mul_2_FpMantRNE_48U_24U_else_and_tmp);
  assign or_235_nl = (~ or_tmp_216) | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign mux_69_nl = MUX_s_1_2_2((or_235_nl), or_tmp_211, mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st);
  assign or_830_nl = (~((FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2
      & mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm) | FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm))
      | (mux_69_nl);
  assign mux_70_nl = MUX_s_1_2_2((or_830_nl), (mux_68_nl), nor_20_cse);
  assign mux_71_nl = MUX_s_1_2_2((mux_70_nl), (or_227_nl), IsNaN_8U_23U_1_land_2_lpi_1_dfm_6);
  assign nor_263_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (mux_71_nl));
  assign nor_268_nl = ~(FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign and_342_nl = mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2
      & FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3
      & (~ FpMul_8U_23U_lor_7_lpi_1_dfm_st_4) & mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign mux_72_nl = MUX_s_1_2_2((and_342_nl), (nor_268_nl), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2);
  assign nand_20_nl = ~((nor_267_cse | mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2)
      & (mux_72_nl));
  assign mux_73_nl = MUX_s_1_2_2((nand_20_nl), IsNaN_8U_23U_land_2_lpi_1_dfm_st_5,
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7);
  assign nor_266_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_8 | mul_mul_land_2_lpi_1_dfm_st_5 | (mux_73_nl));
  assign mux_74_nl = MUX_s_1_2_2((nor_266_nl), (nor_263_nl), or_74_cse);
  assign nor_260_nl = ~((~ (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_2_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | nand_45_cse);
  assign nor_261_nl = ~((~ mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3
      | nand_45_cse);
  assign mux_75_nl = MUX_s_1_2_2((nor_261_nl), (nor_260_nl), nor_20_cse);
  assign nor_262_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 | (~(mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2)));
  assign mux_76_nl = MUX_s_1_2_2((nor_262_nl), (mux_75_nl), or_74_cse);
  assign or_254_nl = nor_264_cse | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_7
      | mul_mul_land_2_lpi_1_dfm_5;
  assign or_255_nl = (~ FpMul_8U_23U_lor_7_lpi_1_dfm_6) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign mux_77_nl = MUX_s_1_2_2((or_255_nl), (or_254_nl), mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_78_nl = MUX_s_1_2_2((mux_77_nl), or_tmp_235, mul_mul_2_FpMantRNE_48U_24U_else_and_tmp);
  assign or_258_nl = (~ or_tmp_216) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_7
      | mul_mul_land_2_lpi_1_dfm_5;
  assign mux_79_nl = MUX_s_1_2_2((or_258_nl), or_tmp_235, mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st);
  assign mux_80_nl = MUX_s_1_2_2((mux_79_nl), (mux_78_nl), nor_20_cse);
  assign nor_255_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (mux_80_nl));
  assign nor_257_nl = ~((~(nor_267_cse | mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2))
      | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_8 | mul_mul_land_2_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_7
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign mux_81_nl = MUX_s_1_2_2((nor_257_nl), (nor_255_nl), or_74_cse);
  assign nor_253_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | nand_45_cse);
  assign nor_254_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 | (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign mux_82_nl = MUX_s_1_2_2((nor_254_nl), (nor_253_nl), or_74_cse);
  assign or_270_nl = or_tmp_252 | or_tmp_167;
  assign mux_84_nl = MUX_s_1_2_2(mux_tmp_78, or_tmp_256, or_tmp_252);
  assign mux_85_nl = MUX_s_1_2_2((mux_84_nl), (or_270_nl), FpMul_8U_23U_lor_7_lpi_1_dfm_st_4);
  assign nor_238_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_2_lpi_1_dfm_7
      | mul_mul_land_2_lpi_1_dfm_5);
  assign nor_240_nl = ~(nor_241_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_2_lpi_1_dfm_7
      | mul_mul_land_2_lpi_1_dfm_5);
  assign nor_242_nl = ~((FpMul_8U_23U_p_mant_p1_2_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5);
  assign mux_90_nl = MUX_s_1_2_2((nor_242_nl), (nor_240_nl), nor_49_cse);
  assign nand_22_nl = ~(mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_90_nl));
  assign or_292_nl = (~ FpMul_8U_23U_FpMul_8U_23U_and_12_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5;
  assign mux_91_nl = MUX_s_1_2_2((or_292_nl), (nand_22_nl), nor_20_cse);
  assign nor_239_nl = ~(FpMul_8U_23U_lor_7_lpi_1_dfm_6 | (mux_91_nl));
  assign mux_92_nl = MUX_s_1_2_2((nor_239_nl), (nor_238_nl), IsNaN_8U_23U_1_land_2_lpi_1_dfm_6);
  assign and_340_nl = (~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | (~ main_stage_v_2))) & (mux_92_nl);
  assign nor_243_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_8 | mul_mul_land_2_lpi_1_dfm_st_5 | (~((~(nor_245_cse
      | FpMul_8U_23U_lor_7_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2)))
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_7)));
  assign mux_93_nl = MUX_s_1_2_2((nor_243_nl), (and_340_nl), or_74_cse);
  assign nor_232_nl = ~(nor_241_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | FpMul_8U_23U_lor_7_lpi_1_dfm_6 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5);
  assign nor_234_nl = ~((FpMul_8U_23U_p_mant_p1_2_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_2_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_7_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5);
  assign mux_95_nl = MUX_s_1_2_2((nor_234_nl), (nor_232_nl), nor_49_cse);
  assign and_339_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_95_nl);
  assign nor_235_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_12_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_2_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_7_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5);
  assign mux_96_nl = MUX_s_1_2_2((nor_235_nl), (and_339_nl), nor_20_cse);
  assign nor_236_nl = ~(nor_245_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5
      | mul_mul_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_8 | mul_mul_land_2_lpi_1_dfm_st_5
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 | FpMul_8U_23U_lor_7_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2));
  assign mux_97_nl = MUX_s_1_2_2((nor_236_nl), (mux_96_nl), or_74_cse);
  assign or_307_nl = IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 | IsNaN_8U_23U_land_3_lpi_1_dfm_7
      | mul_mul_land_3_lpi_1_dfm_5;
  assign or_310_nl = nor_227_cse | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign or_311_nl = (~ FpMul_8U_23U_lor_8_lpi_1_dfm_6) | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3
      | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign mux_98_nl = MUX_s_1_2_2((or_311_nl), (or_310_nl), mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_99_nl = MUX_s_1_2_2((mux_98_nl), or_tmp_291, mul_mul_3_FpMantRNE_48U_24U_else_and_tmp);
  assign or_315_nl = (~ or_tmp_296) | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign mux_100_nl = MUX_s_1_2_2((or_315_nl), or_tmp_291, mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st);
  assign or_829_nl = (~((FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2
      & mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm) | FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm))
      | (mux_100_nl);
  assign mux_101_nl = MUX_s_1_2_2((or_829_nl), (mux_99_nl), nor_20_cse);
  assign mux_102_nl = MUX_s_1_2_2((mux_101_nl), (or_307_nl), IsNaN_8U_23U_1_land_3_lpi_1_dfm_6);
  assign nor_226_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (mux_102_nl));
  assign nor_231_nl = ~(FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign and_338_nl = mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2
      & FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3
      & (~ FpMul_8U_23U_lor_8_lpi_1_dfm_st_4) & mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign mux_103_nl = MUX_s_1_2_2((and_338_nl), (nor_231_nl), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2);
  assign nand_27_nl = ~((nor_230_cse | mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2)
      & (mux_103_nl));
  assign mux_104_nl = MUX_s_1_2_2((nand_27_nl), IsNaN_8U_23U_land_3_lpi_1_dfm_st_5,
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7);
  assign nor_229_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_8 | mul_mul_land_3_lpi_1_dfm_st_5 | (mux_104_nl));
  assign mux_105_nl = MUX_s_1_2_2((nor_229_nl), (nor_226_nl), or_74_cse);
  assign nor_223_nl = ~((~ (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_3_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | nand_42_cse);
  assign nor_224_nl = ~((~ mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3
      | nand_42_cse);
  assign mux_106_nl = MUX_s_1_2_2((nor_224_nl), (nor_223_nl), nor_20_cse);
  assign nor_225_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 | (~(mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2)));
  assign mux_107_nl = MUX_s_1_2_2((nor_225_nl), (mux_106_nl), or_74_cse);
  assign or_334_nl = nor_227_cse | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_7
      | mul_mul_land_3_lpi_1_dfm_5;
  assign or_335_nl = (~ FpMul_8U_23U_lor_8_lpi_1_dfm_6) | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign mux_108_nl = MUX_s_1_2_2((or_335_nl), (or_334_nl), mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_109_nl = MUX_s_1_2_2((mux_108_nl), or_tmp_315, mul_mul_3_FpMantRNE_48U_24U_else_and_tmp);
  assign or_338_nl = (~ or_tmp_296) | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_7
      | mul_mul_land_3_lpi_1_dfm_5;
  assign mux_110_nl = MUX_s_1_2_2((or_338_nl), or_tmp_315, mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st);
  assign mux_111_nl = MUX_s_1_2_2((mux_110_nl), (mux_109_nl), nor_20_cse);
  assign nor_218_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (mux_111_nl));
  assign nor_220_nl = ~((~(nor_230_cse | mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2))
      | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_8 | mul_mul_land_3_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_7
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign mux_112_nl = MUX_s_1_2_2((nor_220_nl), (nor_218_nl), or_74_cse);
  assign nor_216_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | nand_42_cse);
  assign nor_217_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 | (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign mux_113_nl = MUX_s_1_2_2((nor_217_nl), (nor_216_nl), or_74_cse);
  assign or_350_nl = or_tmp_332 | or_tmp_167;
  assign mux_115_nl = MUX_s_1_2_2(mux_tmp_109, or_tmp_336, or_tmp_332);
  assign mux_116_nl = MUX_s_1_2_2((mux_115_nl), (or_350_nl), FpMul_8U_23U_lor_8_lpi_1_dfm_st_4);
  assign nor_201_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_3_lpi_1_dfm_7
      | mul_mul_land_3_lpi_1_dfm_5);
  assign nor_203_nl = ~(nor_204_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_3_lpi_1_dfm_7
      | mul_mul_land_3_lpi_1_dfm_5);
  assign nor_205_nl = ~((FpMul_8U_23U_p_mant_p1_3_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5);
  assign mux_121_nl = MUX_s_1_2_2((nor_205_nl), (nor_203_nl), nor_68_cse);
  assign nand_29_nl = ~(mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_121_nl));
  assign or_372_nl = (~ FpMul_8U_23U_FpMul_8U_23U_and_13_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5;
  assign mux_122_nl = MUX_s_1_2_2((or_372_nl), (nand_29_nl), nor_20_cse);
  assign nor_202_nl = ~(FpMul_8U_23U_lor_8_lpi_1_dfm_6 | (mux_122_nl));
  assign mux_123_nl = MUX_s_1_2_2((nor_202_nl), (nor_201_nl), IsNaN_8U_23U_1_land_3_lpi_1_dfm_6);
  assign and_336_nl = (~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | (~ main_stage_v_2))) & (mux_123_nl);
  assign nor_206_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_8 | mul_mul_land_3_lpi_1_dfm_st_5 | (~((~(nor_208_cse
      | FpMul_8U_23U_lor_8_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2)))
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_7)));
  assign mux_124_nl = MUX_s_1_2_2((nor_206_nl), (and_336_nl), or_74_cse);
  assign nor_195_nl = ~(nor_204_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | FpMul_8U_23U_lor_8_lpi_1_dfm_6 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6
      | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5);
  assign nor_197_nl = ~((FpMul_8U_23U_p_mant_p1_3_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_3_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_8_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5);
  assign mux_126_nl = MUX_s_1_2_2((nor_197_nl), (nor_195_nl), nor_68_cse);
  assign and_335_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_126_nl);
  assign nor_198_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_13_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_3_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_8_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5);
  assign mux_127_nl = MUX_s_1_2_2((nor_198_nl), (and_335_nl), nor_20_cse);
  assign nor_199_nl = ~(nor_208_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5
      | mul_mul_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_8 | mul_mul_land_3_lpi_1_dfm_st_5
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 | FpMul_8U_23U_lor_8_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2));
  assign mux_128_nl = MUX_s_1_2_2((nor_199_nl), (mux_127_nl), or_74_cse);
  assign or_387_nl = IsNaN_8U_23U_land_lpi_1_dfm_st_4 | IsNaN_8U_23U_land_lpi_1_dfm_7
      | mul_mul_land_lpi_1_dfm_5;
  assign or_390_nl = nor_190_cse | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign or_391_nl = (~ FpMul_8U_23U_lor_1_lpi_1_dfm_6) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign mux_129_nl = MUX_s_1_2_2((or_391_nl), (or_390_nl), mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_130_nl = MUX_s_1_2_2((mux_129_nl), or_tmp_371, mul_mul_4_FpMantRNE_48U_24U_else_and_tmp);
  assign or_395_nl = (~ or_tmp_376) | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign mux_131_nl = MUX_s_1_2_2((or_395_nl), or_tmp_371, mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st);
  assign or_828_nl = (~((FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2
      & mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm) | FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm))
      | (mux_131_nl);
  assign mux_132_nl = MUX_s_1_2_2((or_828_nl), (mux_130_nl), nor_20_cse);
  assign mux_133_nl = MUX_s_1_2_2((mux_132_nl), (or_387_nl), IsNaN_8U_23U_1_land_lpi_1_dfm_6);
  assign nor_189_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (mux_133_nl));
  assign nor_194_nl = ~(FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign and_334_nl = mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2
      & FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3
      & (~ FpMul_8U_23U_lor_1_lpi_1_dfm_st_4) & mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign mux_134_nl = MUX_s_1_2_2((and_334_nl), (nor_194_nl), FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2);
  assign nand_34_nl = ~((nor_193_cse | mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2)
      & (mux_134_nl));
  assign mux_135_nl = MUX_s_1_2_2((nand_34_nl), IsNaN_8U_23U_land_lpi_1_dfm_st_5,
      IsNaN_8U_23U_1_land_lpi_1_dfm_7);
  assign nor_192_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_8 | mul_mul_land_lpi_1_dfm_st_5 | (mux_135_nl));
  assign mux_136_nl = MUX_s_1_2_2((nor_192_nl), (nor_189_nl), or_74_cse);
  assign nor_186_nl = ~((~ (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | not_tmp_121);
  assign nor_187_nl = ~((~ mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm)
      | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4 | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3
      | not_tmp_121);
  assign mux_137_nl = MUX_s_1_2_2((nor_187_nl), (nor_186_nl), nor_20_cse);
  assign nor_188_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_lpi_1_dfm_st_5
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | (~(mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4
      & mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2)));
  assign mux_138_nl = MUX_s_1_2_2((nor_188_nl), (mux_137_nl), or_74_cse);
  assign or_414_nl = nor_190_cse | IsNaN_8U_23U_1_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_7
      | mul_mul_land_lpi_1_dfm_5;
  assign or_415_nl = (~ FpMul_8U_23U_lor_1_lpi_1_dfm_6) | IsNaN_8U_23U_1_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign mux_139_nl = MUX_s_1_2_2((or_415_nl), (or_414_nl), mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2);
  assign mux_140_nl = MUX_s_1_2_2((mux_139_nl), or_tmp_395, mul_mul_4_FpMantRNE_48U_24U_else_and_tmp);
  assign or_418_nl = (~ or_tmp_376) | IsNaN_8U_23U_1_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_7
      | mul_mul_land_lpi_1_dfm_5;
  assign mux_141_nl = MUX_s_1_2_2((or_418_nl), or_tmp_395, mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st);
  assign mux_142_nl = MUX_s_1_2_2((mux_141_nl), (mux_140_nl), nor_20_cse);
  assign nor_181_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | (~ main_stage_v_2) | (mux_142_nl));
  assign nor_183_nl = ~((~(nor_193_cse | mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2))
      | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_8 | mul_mul_land_lpi_1_dfm_st_5 | IsNaN_8U_23U_1_land_lpi_1_dfm_7
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4));
  assign mux_143_nl = MUX_s_1_2_2((nor_183_nl), (nor_181_nl), or_74_cse);
  assign or_429_nl = (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | or_tmp_411;
  assign mux_146_nl = MUX_s_1_2_2(mux_tmp_140, or_tmp_415, or_430_cse);
  assign or_424_nl = (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  assign mux_147_nl = MUX_s_1_2_2((mux_146_nl), (or_429_nl), or_424_nl);
  assign or_436_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | or_tmp_411;
  assign mux_148_nl = MUX_s_1_2_2(mux_tmp_140, or_tmp_415, FpMul_8U_23U_lor_1_lpi_1_dfm_st_3);
  assign mux_149_nl = MUX_s_1_2_2((mux_148_nl), (or_436_nl), FpMul_8U_23U_lor_1_lpi_1_dfm_st_4);
  assign nor_167_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_lpi_1_dfm_7
      | mul_mul_land_lpi_1_dfm_5);
  assign nor_169_nl = ~(nor_170_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | IsNaN_8U_23U_land_lpi_1_dfm_7
      | mul_mul_land_lpi_1_dfm_5);
  assign nor_171_nl = ~((FpMul_8U_23U_p_mant_p1_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5);
  assign mux_153_nl = MUX_s_1_2_2((nor_171_nl), (nor_169_nl), nor_86_cse);
  assign nand_36_nl = ~(mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_153_nl));
  assign or_453_nl = (~ FpMul_8U_23U_FpMul_8U_23U_and_14_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5;
  assign mux_154_nl = MUX_s_1_2_2((or_453_nl), (nand_36_nl), nor_20_cse);
  assign nor_168_nl = ~(FpMul_8U_23U_lor_1_lpi_1_dfm_6 | (mux_154_nl));
  assign mux_155_nl = MUX_s_1_2_2((nor_168_nl), (nor_167_nl), IsNaN_8U_23U_1_land_lpi_1_dfm_6);
  assign and_332_nl = (~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | (~ main_stage_v_2))) & (mux_155_nl);
  assign nor_172_nl = ~((~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5 | mul_mul_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_8 | mul_mul_land_lpi_1_dfm_st_5 | (~((~(nor_174_cse
      | FpMul_8U_23U_lor_1_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2)))
      | IsNaN_8U_23U_1_land_lpi_1_dfm_7)));
  assign mux_156_nl = MUX_s_1_2_2((nor_172_nl), (and_332_nl), or_74_cse);
  assign nor_161_nl = ~(nor_170_cse | io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | FpMul_8U_23U_lor_1_lpi_1_dfm_6 | IsNaN_8U_23U_1_land_lpi_1_dfm_6
      | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5);
  assign nor_163_nl = ~((FpMul_8U_23U_p_mant_p1_sva[47]) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_1_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5);
  assign mux_157_nl = MUX_s_1_2_2((nor_163_nl), (nor_161_nl), nor_86_cse);
  assign and_331_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_157_nl);
  assign nor_164_nl = ~((~ FpMul_8U_23U_FpMul_8U_23U_and_14_itm) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_lpi_1_dfm_st_4 | (~ main_stage_v_2) | FpMul_8U_23U_lor_1_lpi_1_dfm_6
      | IsNaN_8U_23U_1_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5);
  assign mux_158_nl = MUX_s_1_2_2((nor_164_nl), (and_331_nl), nor_20_cse);
  assign nor_165_nl = ~(nor_174_cse | (~ main_stage_v_3) | io_read_cfg_mul_bypass_rsc_svs_5
      | mul_mul_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_8 | mul_mul_land_lpi_1_dfm_st_5
      | IsNaN_8U_23U_1_land_lpi_1_dfm_7 | FpMul_8U_23U_lor_1_lpi_1_dfm_7 | (~ FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2));
  assign mux_159_nl = MUX_s_1_2_2((nor_165_nl), (mux_158_nl), or_74_cse);
  assign or_511_nl = (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47]) | mul_mul_land_1_lpi_1_dfm_st_4
      | or_tmp_167;
  assign nor_144_nl = ~((~ (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_land_1_lpi_1_dfm_st_4
      | or_tmp_167);
  assign mux_184_nl = MUX_s_1_2_2((nor_144_nl), (or_511_nl), mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign or_509_nl = (cfg_precision!=2'b10) | (~ mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign mux_185_nl = MUX_s_1_2_2((mux_184_nl), mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_509_nl);
  assign or_515_nl = (~ (mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  assign mux_186_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_1_sva[47])), (or_515_nl),
      nor_31_cse);
  assign and_39_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_186_nl);
  assign nor_100_nl = ~(nor_143_cse | (cfg_precision!=2'b10) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_1_lpi_1_dfm_st_4 | (~ main_stage_v_2));
  assign mux_187_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_itm, (and_39_nl),
      nor_100_nl);
  assign or_519_nl = (~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_mul_land_2_lpi_1_dfm_st_4 | or_tmp_167;
  assign nor_142_nl = ~((~ mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (~ (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_mul_land_2_lpi_1_dfm_st_4 | or_tmp_167);
  assign mux_188_nl = MUX_s_1_2_2((nor_142_nl), (or_519_nl), mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_189_nl = MUX_s_1_2_2((mux_188_nl), mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_27_cse);
  assign or_523_nl = (~ (mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  assign mux_190_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_2_sva[47])), (or_523_nl),
      nor_49_cse);
  assign and_40_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_190_nl);
  assign nor_102_nl = ~(nor_143_cse | (cfg_precision!=2'b10) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_2_lpi_1_dfm_st_4 | (~ main_stage_v_2));
  assign mux_191_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_12_itm, (and_40_nl),
      nor_102_nl);
  assign or_527_nl = (~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | mul_mul_land_3_lpi_1_dfm_st_4 | or_tmp_167;
  assign nor_140_nl = ~((~ mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (~ (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | mul_mul_land_3_lpi_1_dfm_st_4 | or_tmp_167);
  assign mux_192_nl = MUX_s_1_2_2((nor_140_nl), (or_527_nl), mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_193_nl = MUX_s_1_2_2((mux_192_nl), mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_27_cse);
  assign or_531_nl = (~ (mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47])) | mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  assign mux_194_nl = MUX_s_1_2_2((~ (FpMul_8U_23U_p_mant_p1_3_sva[47])), (or_531_nl),
      nor_68_cse);
  assign and_41_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2
      & (mux_194_nl);
  assign nor_104_nl = ~(nor_143_cse | (cfg_precision!=2'b10) | io_read_cfg_mul_bypass_rsc_svs_st_4
      | mul_mul_land_3_lpi_1_dfm_st_4 | (~ main_stage_v_2));
  assign mux_195_nl = MUX_s_1_2_2(FpMul_8U_23U_FpMul_8U_23U_and_13_itm, (and_41_nl),
      nor_104_nl);
  assign or_535_nl = (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47])
      | or_tmp_411;
  assign nor_342_nl = ~((~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (~ (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))
      | or_tmp_411);
  assign mux_196_nl = MUX_s_1_2_2((nor_342_nl), (or_535_nl), mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm);
  assign mux_197_nl = MUX_s_1_2_2((mux_196_nl), mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm,
      or_27_cse);
  assign nor_107_nl = ~((FpMul_8U_23U_p_mant_p1_sva[47]) | (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2));
  assign mux_198_nl = MUX_s_1_2_2(and_tmp_5, or_tmp_517, nor_107_nl);
  assign and_328_nl = (mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 | (~
      (mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47]))) & mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign mux_199_nl = MUX_s_1_2_2(and_tmp_5, or_tmp_517, and_328_nl);
  assign mux_200_nl = MUX_s_1_2_2((mux_199_nl), (mux_198_nl), or_430_cse);
  assign mux_201_nl = MUX_s_1_2_2((mux_200_nl), FpMul_8U_23U_FpMul_8U_23U_and_14_itm,
      or_27_cse);
  assign FpMul_8U_23U_oelse_1_mux_20_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_6_lpi_1_dfm_6,
      FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0, and_18_tmp);
  assign nor_136_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_1_lpi_1_dfm_st_1
      | IsNaN_8U_23U_land_1_lpi_1_dfm_4 | mul_mul_land_1_lpi_1_dfm_2);
  assign nor_137_nl = ~(((~ IsNaN_8U_23U_1_nor_tmp) & (else_mux_tmp_30_23==8'b11111111))
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_1_lpi_1_dfm_st_1 | IsNaN_8U_23U_land_1_lpi_1_dfm_4
      | mul_mul_land_1_lpi_1_dfm_2);
  assign or_540_nl = (cfg_precision!=2'b10) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_1;
  assign mux_202_nl = MUX_s_1_2_2((nor_137_nl), (nor_136_nl), or_540_nl);
  assign nor_138_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_1_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_land_1_lpi_1_dfm_7 | mul_mul_land_1_lpi_1_dfm_5);
  assign mux_203_nl = MUX_s_1_2_2((nor_138_nl), (mux_202_nl), and_18_tmp);
  assign mul_mul_1_FpMul_8U_23U_xor_nl = (MulIn_data_sva_1[31]) ^ (else_MulOp_data_0_lpi_1_dfm_mx1[31]);
  assign nor_134_nl = ~(mul_mul_land_1_lpi_1_dfm_2 | io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_135_nl = ~((~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mul_mul_land_1_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2));
  assign mux_207_nl = MUX_s_1_2_2((nor_135_nl), (nor_134_nl), and_18_tmp);
  assign FpMul_8U_23U_oelse_1_mux_21_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_7_lpi_1_dfm_6,
      FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0, and_18_tmp);
  assign nor_131_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_2_lpi_1_dfm_st_1
      | IsNaN_8U_23U_land_2_lpi_1_dfm_4 | mul_mul_land_2_lpi_1_dfm_2);
  assign nor_132_nl = ~(((~ IsNaN_8U_23U_1_nor_1_tmp) & (else_mux_1_tmp_30_23==8'b11111111))
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_2_lpi_1_dfm_st_1 | IsNaN_8U_23U_land_2_lpi_1_dfm_4
      | mul_mul_land_2_lpi_1_dfm_2);
  assign or_551_nl = (cfg_precision!=2'b10) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_1;
  assign mux_208_nl = MUX_s_1_2_2((nor_132_nl), (nor_131_nl), or_551_nl);
  assign nor_133_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_2_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_land_2_lpi_1_dfm_7 | mul_mul_land_2_lpi_1_dfm_5);
  assign mux_209_nl = MUX_s_1_2_2((nor_133_nl), (mux_208_nl), and_18_tmp);
  assign mul_mul_2_FpMul_8U_23U_xor_nl = (MulIn_data_sva_1[63]) ^ (else_MulOp_data_1_lpi_1_dfm_mx1[31]);
  assign nor_129_nl = ~(mul_mul_land_2_lpi_1_dfm_2 | io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_130_nl = ~((~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mul_mul_land_2_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2));
  assign mux_213_nl = MUX_s_1_2_2((nor_130_nl), (nor_129_nl), and_18_tmp);
  assign FpMul_8U_23U_oelse_1_mux_22_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_8_lpi_1_dfm_6,
      FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0, and_18_tmp);
  assign nor_126_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_3_lpi_1_dfm_st_1
      | IsNaN_8U_23U_land_3_lpi_1_dfm_4 | mul_mul_land_3_lpi_1_dfm_2);
  assign nor_127_nl = ~(((~ IsNaN_8U_23U_1_nor_2_tmp) & (else_mux_2_tmp_30_23==8'b11111111))
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_3_lpi_1_dfm_st_1 | IsNaN_8U_23U_land_3_lpi_1_dfm_4
      | mul_mul_land_3_lpi_1_dfm_2);
  assign or_561_nl = (cfg_precision!=2'b10) | IsNaN_8U_23U_land_3_lpi_1_dfm_st_1;
  assign mux_214_nl = MUX_s_1_2_2((nor_127_nl), (nor_126_nl), or_561_nl);
  assign nor_128_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_3_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_land_3_lpi_1_dfm_7 | mul_mul_land_3_lpi_1_dfm_5);
  assign mux_215_nl = MUX_s_1_2_2((nor_128_nl), (mux_214_nl), and_18_tmp);
  assign mul_mul_3_FpMul_8U_23U_xor_nl = (MulIn_data_sva_1[95]) ^ (else_MulOp_data_2_lpi_1_dfm_mx1[31]);
  assign nor_124_nl = ~(mul_mul_land_3_lpi_1_dfm_2 | io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_125_nl = ~((~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mul_mul_land_3_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2));
  assign mux_219_nl = MUX_s_1_2_2((nor_125_nl), (nor_124_nl), and_18_tmp);
  assign FpMul_8U_23U_oelse_1_mux_23_nl = MUX_s_1_2_2(FpMul_8U_23U_lor_1_lpi_1_dfm_6,
      FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0, and_18_tmp);
  assign nor_121_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_lpi_1_dfm_st_1
      | IsNaN_8U_23U_land_lpi_1_dfm_4 | mul_mul_land_lpi_1_dfm_2);
  assign nor_122_nl = ~(((~ IsNaN_8U_23U_1_nor_3_tmp) & (else_mux_3_tmp_30_23==8'b11111111))
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_land_lpi_1_dfm_st_1 | IsNaN_8U_23U_land_lpi_1_dfm_4
      | mul_mul_land_lpi_1_dfm_2);
  assign or_571_nl = (cfg_precision!=2'b10) | IsNaN_8U_23U_land_lpi_1_dfm_st_1;
  assign mux_220_nl = MUX_s_1_2_2((nor_122_nl), (nor_121_nl), or_571_nl);
  assign nor_123_nl = ~(io_read_cfg_mul_bypass_rsc_svs_st_4 | mul_mul_land_lpi_1_dfm_st_4
      | (~ main_stage_v_2) | (~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | IsNaN_8U_23U_1_land_lpi_1_dfm_6 | IsNaN_8U_23U_land_lpi_1_dfm_7 | mul_mul_land_lpi_1_dfm_5);
  assign mux_221_nl = MUX_s_1_2_2((nor_123_nl), (mux_220_nl), and_18_tmp);
  assign mul_mul_4_FpMul_8U_23U_xor_nl = (MulIn_data_sva_1[127]) ^ (else_MulOp_data_3_lpi_1_dfm_mx1[31]);
  assign nor_119_nl = ~(mul_mul_land_lpi_1_dfm_2 | io_read_cfg_mul_bypass_rsc_svs_st_1);
  assign nor_120_nl = ~((~ reg_chn_mul_out_rsci_ld_core_psct_cse) | chn_mul_out_rsci_bawt
      | mul_mul_land_lpi_1_dfm_5 | io_read_cfg_mul_bypass_rsc_svs_st_4 | (~ main_stage_v_2));
  assign mux_225_nl = MUX_s_1_2_2((nor_120_nl), (nor_119_nl), and_18_tmp);
  assign nor_159_nl = ~(or_tmp_1 | nor_118_cse);
  assign mux_161_nl = MUX_s_1_2_2((nor_159_nl), or_tmp_12, FpMul_8U_23U_lor_6_lpi_1_dfm_st);
  assign or_473_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st | (~ or_tmp_1);
  assign mux_162_nl = MUX_s_1_2_2((or_473_nl), (mux_161_nl), mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign or_474_nl = (~ mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1) | mul_mul_land_1_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | IsZero_8U_23U_land_1_lpi_1_dfm_4 |
      mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  assign mux_163_nl = MUX_s_1_2_2((or_474_nl), (mux_162_nl), mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs);
  assign mux_164_nl = MUX_s_1_2_2((mux_163_nl), or_469_cse, or_468_cse);
  assign nor_157_nl = ~(or_tmp_15 | nor_117_cse);
  assign mux_169_nl = MUX_s_1_2_2((nor_157_nl), or_tmp_26, FpMul_8U_23U_lor_7_lpi_1_dfm_st);
  assign or_486_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st | (~ or_tmp_15);
  assign mux_170_nl = MUX_s_1_2_2((or_486_nl), (mux_169_nl), mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign or_487_nl = (~ mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1) | mul_mul_land_2_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | IsZero_8U_23U_land_2_lpi_1_dfm_4 |
      mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  assign mux_171_nl = MUX_s_1_2_2((or_487_nl), (mux_170_nl), mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs);
  assign mux_172_nl = MUX_s_1_2_2((mux_171_nl), or_482_cse, or_468_cse);
  assign nor_155_nl = ~(or_tmp_29 | nor_116_cse);
  assign mux_174_nl = MUX_s_1_2_2((nor_155_nl), or_tmp_40, FpMul_8U_23U_lor_8_lpi_1_dfm_st);
  assign or_494_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st | (~ or_tmp_29);
  assign mux_175_nl = MUX_s_1_2_2((or_494_nl), (mux_174_nl), mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign or_495_nl = (~ mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1) | mul_mul_land_3_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | IsZero_8U_23U_land_3_lpi_1_dfm_4 |
      mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  assign mux_176_nl = MUX_s_1_2_2((or_495_nl), (mux_175_nl), mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs);
  assign mux_177_nl = MUX_s_1_2_2((mux_176_nl), or_490_cse, or_468_cse);
  assign or_498_nl = (~ mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs)
      | FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  assign nor_153_nl = ~(or_tmp_46 | nor_115_cse);
  assign mux_179_nl = MUX_s_1_2_2((nor_153_nl), or_tmp_51, FpMul_8U_23U_lor_1_lpi_1_dfm_st);
  assign or_502_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st | (~ or_tmp_46);
  assign mux_180_nl = MUX_s_1_2_2((or_502_nl), (mux_179_nl), mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1);
  assign or_503_nl = (~ mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1) | mul_mul_land_lpi_1_dfm_st_1
      | io_read_cfg_mul_bypass_rsc_svs_st_1 | mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1
      | IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp | IsZero_8U_23U_land_lpi_1_dfm_4;
  assign mux_181_nl = MUX_s_1_2_2((or_503_nl), (mux_180_nl), mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs);
  assign mux_182_nl = MUX_s_1_2_2((mux_181_nl), (or_498_nl), or_468_cse);

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [21:0] MUX1HOT_v_22_3_2;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [2:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    MUX1HOT_v_22_3_2 = result;
  end
  endfunction


  function [22:0] MUX1HOT_v_23_3_2;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [2:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    MUX1HOT_v_23_3_2 = result;
  end
  endfunction


  function [22:0] MUX1HOT_v_23_4_2;
    input [22:0] input_3;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [3:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    result = result | ( input_3 & {23{sel[3]}});
    MUX1HOT_v_23_4_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [45:0] MUX_v_46_2_2;
    input [45:0] input_0;
    input [45:0] input_1;
    input [0:0] sel;
    reg [45:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_46_2_2 = result;
  end
  endfunction


  function [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function [22:0] signext_23_1;
    input [0:0] vector;
  begin
    signext_23_1= {{22{vector[0]}}, vector};
  end
  endfunction


  function  [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function  [64:0] conv_s2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_s2s_64_65 = {vector[63], vector};
  end
  endfunction


  function  [63:0] conv_s2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_s2u_64_64 = vector;
  end
  endfunction


  function  [64:0] conv_u2s_1_65 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_65 = {{64{1'b0}}, vector};
  end
  endfunction


  function  [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function  [9:0] conv_u2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [22:0] conv_u2u_1_23 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction


  function  [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function  [47:0] conv_u2u_48_48 ;
    input [47:0]  vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu_core
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu_core (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz,
      chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, cfg_alu_bypass_rsc_triosy_lz,
      cfg_alu_src_rsc_triosy_lz, cfg_alu_op_rsc_triosy_lz, cfg_alu_algo_rsc_triosy_lz,
      cfg_precision, chn_alu_out_rsc_z, chn_alu_out_rsc_vz, chn_alu_out_rsc_lz, chn_alu_in_rsci_oswt,
      chn_alu_in_rsci_oswt_unreg, chn_alu_op_rsci_oswt, chn_alu_op_rsci_oswt_unreg,
      cfg_alu_bypass_rsci_d, cfg_alu_src_rsci_d, cfg_alu_op_rsci_d, cfg_alu_algo_rsci_d,
      chn_alu_out_rsci_oswt, chn_alu_out_rsci_oswt_unreg, cfg_alu_bypass_rsc_triosy_obj_oswt,
      cfg_alu_src_rsc_triosy_obj_oswt, cfg_alu_op_rsc_triosy_obj_oswt, cfg_alu_algo_rsc_triosy_obj_oswt,
      cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_alu_in_rsc_z;
  input chn_alu_in_rsc_vz;
  output chn_alu_in_rsc_lz;
  input [127:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  output cfg_alu_bypass_rsc_triosy_lz;
  output cfg_alu_src_rsc_triosy_lz;
  output cfg_alu_op_rsc_triosy_lz;
  output cfg_alu_algo_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [127:0] chn_alu_out_rsc_z;
  input chn_alu_out_rsc_vz;
  output chn_alu_out_rsc_lz;
  input chn_alu_in_rsci_oswt;
  output chn_alu_in_rsci_oswt_unreg;
  input chn_alu_op_rsci_oswt;
  output chn_alu_op_rsci_oswt_unreg;
  input cfg_alu_bypass_rsci_d;
  input cfg_alu_src_rsci_d;
  input [31:0] cfg_alu_op_rsci_d;
  input [1:0] cfg_alu_algo_rsci_d;
  input chn_alu_out_rsci_oswt;
  output chn_alu_out_rsci_oswt_unreg;
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  input cfg_alu_src_rsc_triosy_obj_oswt;
  input cfg_alu_op_rsc_triosy_obj_oswt;
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  output cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff;


  // Interconnect Declarations
  wire core_wen;
  reg chn_alu_in_rsci_iswt0;
  wire chn_alu_in_rsci_bawt;
  wire chn_alu_in_rsci_wen_comp;
  reg chn_alu_in_rsci_ld_core_psct;
  wire [127:0] chn_alu_in_rsci_d_mxwt;
  wire core_wten;
  reg chn_alu_op_rsci_iswt0;
  wire chn_alu_op_rsci_bawt;
  wire chn_alu_op_rsci_wen_comp;
  reg chn_alu_op_rsci_ld_core_psct;
  wire [127:0] chn_alu_op_rsci_d_mxwt;
  reg chn_alu_out_rsci_iswt0;
  wire chn_alu_out_rsci_bawt;
  wire chn_alu_out_rsci_wen_comp;
  wire cfg_alu_bypass_rsc_triosy_obj_bawt;
  wire cfg_alu_src_rsc_triosy_obj_bawt;
  wire cfg_alu_op_rsc_triosy_obj_bawt;
  wire cfg_alu_algo_rsc_triosy_obj_bawt;
  reg chn_alu_out_rsci_d_127;
  reg [7:0] chn_alu_out_rsci_d_126_119;
  reg [21:0] chn_alu_out_rsci_d_118_97;
  reg chn_alu_out_rsci_d_96;
  reg chn_alu_out_rsci_d_95;
  reg [7:0] chn_alu_out_rsci_d_94_87;
  reg [21:0] chn_alu_out_rsci_d_86_65;
  reg chn_alu_out_rsci_d_64;
  reg chn_alu_out_rsci_d_63;
  reg [7:0] chn_alu_out_rsci_d_62_55;
  reg [21:0] chn_alu_out_rsci_d_54_33;
  reg chn_alu_out_rsci_d_32;
  reg chn_alu_out_rsci_d_31;
  reg [7:0] chn_alu_out_rsci_d_30_23;
  reg [21:0] chn_alu_out_rsci_d_22_1;
  reg chn_alu_out_rsci_d_0;
  wire [1:0] fsm_output;
  wire alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp;
  wire alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp;
  wire alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp;
  wire alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp;
  wire alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
  wire alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
  wire alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
  wire alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  wire IsNaN_8U_23U_3_nor_10_tmp;
  wire IsNaN_8U_23U_3_nor_8_tmp;
  wire IsNaN_8U_23U_3_nor_6_tmp;
  wire IsNaN_8U_23U_3_nor_4_tmp;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_tmp;
  wire or_tmp_9;
  wire mux_tmp_2;
  wire or_tmp_15;
  wire mux_tmp_10;
  wire or_tmp_20;
  wire not_tmp_24;
  wire or_tmp_23;
  wire not_tmp_29;
  wire not_tmp_38;
  wire or_tmp_75;
  wire not_tmp_57;
  wire or_tmp_103;
  wire mux_tmp_53;
  wire or_tmp_218;
  wire or_tmp_224;
  wire or_tmp_251;
  wire or_tmp_261;
  wire or_tmp_269;
  wire or_tmp_280;
  wire or_tmp_293;
  wire or_tmp_305;
  wire or_tmp_309;
  wire or_tmp_312;
  wire or_tmp_315;
  wire or_tmp_347;
  wire not_tmp_152;
  wire mux_tmp_146;
  wire nand_tmp_13;
  wire not_tmp_157;
  wire or_tmp_382;
  wire or_tmp_386;
  wire nor_tmp_74;
  wire or_tmp_395;
  wire mux_tmp_164;
  wire mux_tmp_165;
  wire or_tmp_402;
  wire mux_tmp_171;
  wire or_tmp_409;
  wire mux_tmp_173;
  wire or_tmp_416;
  wire not_tmp_232;
  wire or_tmp_577;
  wire mux_tmp_227;
  wire or_tmp_583;
  wire or_tmp_585;
  wire mux_tmp_237;
  wire nand_tmp_20;
  wire mux_tmp_246;
  wire not_tmp_259;
  wire or_tmp_596;
  wire or_tmp_597;
  wire not_tmp_261;
  wire mux_tmp_265;
  wire mux_tmp_268;
  wire mux_tmp_281;
  wire nor_tmp_126;
  wire and_tmp_35;
  wire mux_tmp_296;
  wire or_dcpl_14;
  wire and_dcpl_28;
  wire and_dcpl_30;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire or_dcpl_20;
  wire and_dcpl_35;
  wire and_dcpl_37;
  wire and_dcpl_40;
  wire or_dcpl_23;
  wire and_dcpl_43;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_53;
  wire and_dcpl_64;
  wire and_dcpl_70;
  wire or_dcpl_46;
  wire or_dcpl_49;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_83;
  wire and_dcpl_89;
  wire and_dcpl_96;
  wire and_dcpl_99;
  wire and_dcpl_108;
  wire or_tmp_657;
  wire mux_tmp_311;
  wire nor_tmp_144;
  wire and_dcpl_127;
  wire or_dcpl_85;
  wire or_dcpl_86;
  wire or_dcpl_89;
  wire or_dcpl_91;
  wire or_dcpl_100;
  wire or_dcpl_109;
  wire or_dcpl_117;
  wire or_dcpl_119;
  wire or_dcpl_121;
  wire or_dcpl_123;
  wire and_dcpl_165;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire or_dcpl_125;
  wire or_dcpl_127;
  wire and_dcpl_175;
  wire and_dcpl_179;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire mux_tmp_323;
  wire and_dcpl_214;
  wire and_dcpl_217;
  wire and_dcpl_219;
  wire and_dcpl_222;
  wire and_dcpl_225;
  wire or_dcpl_154;
  wire and_dcpl_227;
  wire and_dcpl_229;
  wire and_dcpl_231;
  wire and_dcpl_234;
  wire and_dcpl_236;
  wire and_dcpl_239;
  wire and_dcpl_243;
  wire or_tmp_668;
  wire or_tmp_674;
  wire or_tmp_678;
  wire or_tmp_695;
  reg [7:0] FpAdd_8U_23U_qr_2_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_qr_3_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_qr_4_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_qr_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm;
  reg FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2;
  reg alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  reg [7:0] FpAlu_8U_23U_o_30_23_lpi_1_dfm_4;
  reg [21:0] FpAlu_8U_23U_o_22_1_lpi_1_dfm_4;
  reg FpAlu_8U_23U_o_0_lpi_1_dfm_4;
  reg [7:0] AluOut_data_2_30_23_lpi_1_dfm_3;
  reg [21:0] AluOut_data_2_22_1_lpi_1_dfm_3;
  reg AluOut_data_2_0_lpi_1_dfm_3;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  reg FpAdd_8U_23U_and_2_tmp_3;
  reg [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13;
  reg FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  reg FpAdd_8U_23U_and_1_tmp_3;
  reg [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13;
  reg FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  reg FpAdd_8U_23U_and_tmp_2;
  reg [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13;
  reg FpAdd_8U_23U_is_inf_lpi_1_dfm_8;
  reg FpAdd_8U_23U_and_3_tmp_3;
  reg [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_13;
  reg FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6;
  reg FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6;
  reg FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6;
  reg FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  reg IsNaN_8U_23U_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_land_lpi_1_dfm_9;
  reg IsNaN_8U_23U_land_lpi_1_dfm_10;
  reg IsNaN_8U_23U_land_lpi_1_dfm_11;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  reg alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  reg alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  reg FpAlu_8U_23U_equal_tmp_21;
  reg FpAlu_8U_23U_equal_tmp_22;
  reg FpAlu_8U_23U_equal_tmp_23;
  reg FpAlu_8U_23U_equal_tmp_24;
  reg FpAlu_8U_23U_equal_tmp_25;
  reg FpAlu_8U_23U_equal_tmp_26;
  reg FpAlu_8U_23U_nor_dfs_4;
  reg FpAlu_8U_23U_nor_dfs_5;
  reg FpAlu_8U_23U_nor_dfs_6;
  reg FpAlu_8U_23U_equal_tmp_27;
  reg FpAlu_8U_23U_equal_tmp_28;
  reg FpAlu_8U_23U_equal_tmp_29;
  reg FpAlu_8U_23U_equal_tmp_30;
  reg FpAlu_8U_23U_equal_tmp_31;
  reg FpAlu_8U_23U_equal_tmp_32;
  reg FpAlu_8U_23U_equal_tmp_33;
  reg FpAlu_8U_23U_equal_tmp_34;
  reg FpAlu_8U_23U_equal_tmp_35;
  reg alu_loop_op_unequal_tmp_6;
  reg alu_loop_op_unequal_tmp_7;
  reg alu_loop_op_unequal_tmp_8;
  reg FpAlu_8U_23U_o_0_sva_7;
  reg FpAlu_8U_23U_o_0_sva_8;
  reg FpAlu_8U_23U_o_0_sva_9;
  reg AluOut_data_2_0_sva_9;
  reg AluOut_data_2_0_sva_10;
  reg AluOut_data_2_0_sva_11;
  reg AluOut_data_1_0_sva_10;
  reg AluOut_data_1_0_sva_11;
  reg AluOut_data_1_0_sva_12;
  reg AluOut_data_0_0_sva_9;
  reg AluOut_data_0_0_sva_10;
  reg AluOut_data_0_0_sva_11;
  reg [31:0] cfg_alu_op_1_sva_1;
  reg [1:0] cfg_alu_algo_1_sva_2;
  reg [127:0] AluIn_data_sva_127;
  reg [127:0] AluIn_data_sva_128;
  reg io_read_cfg_alu_bypass_rsc_svs_5;
  reg io_read_cfg_alu_bypass_rsc_svs_6;
  reg io_read_cfg_alu_bypass_rsc_svs_7;
  reg io_read_cfg_alu_bypass_rsc_svs_8;
  reg [7:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_6;
  reg [7:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_7;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_6;
  reg [7:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_7;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_6;
  reg [7:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_7;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_qr_lpi_1_dfm_6;
  reg [7:0] FpAdd_8U_23U_qr_lpi_1_dfm_7;
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5;
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5;
  reg [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5;
  reg alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  reg alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  reg AluOut_data_2_31_lpi_1_dfm_6;
  reg AluOut_data_2_31_lpi_1_dfm_7;
  reg cfg_alu_src_1_sva_st;
  reg [1:0] cfg_alu_algo_1_sva_st;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  reg alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  reg alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  reg FpNormalize_8U_49U_if_or_itm;
  reg FpNormalize_8U_49U_if_or_itm_2;
  reg alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st;
  reg alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  reg alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st;
  reg alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm;
  reg FpNormalize_8U_49U_if_or_1_itm;
  reg FpNormalize_8U_49U_if_or_1_itm_2;
  reg alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st;
  reg alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  reg alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  reg alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  reg FpNormalize_8U_49U_if_or_2_itm;
  reg FpNormalize_8U_49U_if_or_2_itm_2;
  reg alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st;
  reg alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  reg alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st;
  reg alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm;
  reg FpNormalize_8U_49U_if_or_3_itm;
  reg FpNormalize_8U_49U_if_or_3_itm_2;
  reg alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st;
  reg alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm;
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm;
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
  reg [1:0] cfg_alu_algo_1_sva_st_20;
  reg IsNaN_8U_23U_4_nor_2_itm_2;
  reg IsNaN_8U_23U_4_nor_3_itm_2;
  reg IsNaN_8U_23U_4_nor_3_itm_3;
  reg FpAlu_8U_23U_mux1h_33_itm_2;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm;
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3;
  reg FpAlu_8U_23U_mux1h_152_itm_2;
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4;
  reg mux_189_itm_3;
  reg mux_189_itm_4;
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4;
  reg FpAlu_8U_23U_and_6_itm_2;
  reg mux_181_itm_3;
  reg mux_181_itm_4;
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4;
  reg FpAlu_8U_23U_and_3_itm_2;
  reg mux_177_itm_3;
  reg mux_177_itm_4;
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2;
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2;
  reg io_read_cfg_alu_bypass_rsc_svs_st_1;
  reg cfg_alu_src_1_sva_st_1;
  reg [1:0] cfg_alu_algo_1_sva_st_22;
  reg io_read_cfg_alu_bypass_rsc_svs_st_5;
  reg [1:0] cfg_alu_algo_1_sva_st_23;
  reg io_read_cfg_alu_bypass_rsc_svs_st_6;
  reg [1:0] cfg_alu_algo_1_sva_st_24;
  reg alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  reg io_read_cfg_alu_bypass_rsc_svs_st_7;
  reg [1:0] cfg_alu_algo_1_sva_st_25;
  reg alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2;
  reg alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  reg alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2;
  reg alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2;
  reg alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  reg alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  reg alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2;
  reg alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  reg alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2;
  reg alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2;
  reg alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  reg [1:0] cfg_alu_algo_1_sva_st_28;
  reg [30:0] else_AluOp_data_0_lpi_1_dfm_2_30_0_1;
  reg [30:0] else_AluOp_data_2_lpi_1_dfm_2_30_0_1;
  reg [30:0] else_AluOp_data_1_lpi_1_dfm_2_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1;
  reg [30:0] FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1;
  reg [30:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1;
  reg [30:0] AluIn_data_sva_3_126_96_1;
  reg [30:0] AluIn_data_sva_3_94_64_1;
  reg [30:0] AluIn_data_sva_3_62_32_1;
  reg [30:0] AluIn_data_sva_3_30_0_1;
  reg [30:0] else_AluOp_data_3_lpi_1_dfm_2_30_0_1;
  wire [8:0] else_mux_3_tmp_31_23;
  wire [8:0] else_mux_2_tmp_31_23;
  wire [8:0] else_mux_1_tmp_31_23;
  wire [8:0] else_mux_tmp_31_23;
  wire and_357_cse;
  wire main_stage_en_1;
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c;
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c;
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c;
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c;
  wire FpAlu_8U_23U_and_12_tmp;
  wire FpAlu_8U_23U_equal_tmp_2_mx0w0;
  wire FpAlu_8U_23U_equal_tmp_1_mx0w0;
  wire alu_loop_op_else_equal_tmp_2;
  wire IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  wire FpAlu_8U_23U_and_38_m1c;
  wire FpAlu_8U_23U_nor_dfs_mx0w0;
  wire IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
  wire FpAlu_8U_23U_and_36_m1c;
  wire IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
  wire FpAlu_8U_23U_and_34_m1c;
  wire IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0;
  wire FpAlu_8U_23U_and_24_m1c;
  wire FpAlu_8U_23U_equal_tmp_mx0w0;
  wire FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0;
  wire IsNaN_8U_23U_2_nor_3_mx0w0;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2;
  wire IsNaN_8U_23U_2_nor_2_mx0w0;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2;
  wire [31:0] else_AluOp_data_3_lpi_1_dfm_mx0;
  wire [31:0] else_AluOp_data_2_lpi_1_dfm_mx0;
  wire [31:0] else_AluOp_data_1_lpi_1_dfm_mx0;
  wire [31:0] else_AluOp_data_0_lpi_1_dfm_mx0;
  wire [30:0] else_AluOp_data_2_lpi_1_dfm_mx3_30_0;
  wire [30:0] else_AluOp_data_0_lpi_1_dfm_mx3_30_0;
  wire and_297_m1c;
  wire chn_alu_out_and_1_cse;
  wire chn_alu_out_and_cse;
  wire chn_alu_out_and_8_cse;
  reg reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse;
  wire nor_6_cse;
  reg reg_chn_alu_out_rsci_ld_core_psct_cse;
  wire FpMantRNE_49U_24U_else_and_cse;
  wire nor_264_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_cse;
  wire FpAdd_8U_23U_if_3_and_cse;
  wire FpAdd_8U_23U_is_addition_and_cse;
  wire nor_269_cse;
  wire nor_236_cse;
  wire alu_loop_bypass_if_and_6_cse;
  wire alu_loop_bypass_if_and_7_cse;
  wire or_963_cse;
  wire AluOut_data_and_5_cse;
  wire nor_202_cse;
  wire or_937_cse;
  wire IsNaN_8U_23U_2_and_cse;
  wire and_486_cse;
  wire nor_5_cse;
  wire and_451_cse;
  wire nor_33_cse;
  wire nor_37_cse;
  wire nor_41_cse;
  wire nor_45_cse;
  wire or_861_cse;
  wire or_867_cse;
  wire or_871_cse;
  wire nor_197_cse;
  wire or_391_cse;
  wire or_381_cse;
  wire and_484_cse;
  wire mux_312_cse;
  wire mux_282_cse;
  wire or_632_cse;
  wire or_28_cse;
  wire FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  wire FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  wire FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  wire FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  wire and_481_cse;
  wire and_501_cse;
  wire nor_177_cse;
  wire nor_71_cse;
  wire and_37_cse;
  wire nor_201_cse;
  wire or_16_cse;
  wire nor_397_cse;
  wire IsZero_8U_23U_1_and_cse;
  wire and_489_cse;
  wire and_524_cse;
  wire and_dcpl_269;
  wire asn_267;
  wire or_997_tmp;
  wire or_996_tmp;
  wire or_998_tmp;
  wire and_167_rgt;
  wire and_dcpl;
  wire and_211_rgt;
  wire and_213_rgt;
  wire and_215_rgt;
  wire and_217_rgt;
  wire and_231_rgt;
  wire and_233_rgt;
  wire and_235_rgt;
  wire and_237_rgt;
  wire and_239_rgt;
  wire and_241_rgt;
  wire and_243_rgt;
  wire and_245_rgt;
  wire and_dcpl_349;
  wire and_293_rgt;
  wire and_328_rgt;
  wire [30:0] AluIn_data_mux1h_7_itm;
  reg [7:0] reg_AluIn_data_sva_4_126_96_itm;
  reg [22:0] reg_AluIn_data_sva_4_126_96_1_itm;
  wire [30:0] AluIn_data_mux1h_9_itm;
  reg [7:0] reg_AluIn_data_sva_4_94_64_itm;
  reg [22:0] reg_AluIn_data_sva_4_94_64_1_itm;
  wire [30:0] AluIn_data_mux1h_11_itm;
  reg [7:0] reg_AluIn_data_sva_4_62_32_itm;
  reg [22:0] reg_AluIn_data_sva_4_62_32_1_itm;
  wire [30:0] AluIn_data_mux1h_13_itm;
  reg [7:0] reg_AluIn_data_sva_4_30_0_itm;
  reg [22:0] reg_AluIn_data_sva_4_30_0_1_itm;
  wire [31:0] alu_loop_op_else_o_mux1h_1_itm;
  reg reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm;
  reg [30:0] reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm;
  wire [31:0] alu_loop_op_else_o_mux1h_3_itm;
  reg reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm;
  reg [30:0] reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm;
  wire [31:0] alu_loop_op_else_o_mux1h_5_itm;
  reg reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm;
  reg [30:0] reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm;
  wire [31:0] alu_loop_op_else_o_mux1h_7_itm;
  reg reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm;
  reg [30:0] reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm;
  wire [48:0] alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_itm;
  wire [48:0] alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_itm;
  wire [48:0] alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_itm;
  wire [48:0] alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm;
  wire mux_34_itm;
  wire mux_109_itm;
  wire mux_143_itm;
  wire mux_337_itm;
  wire FpAdd_8U_23U_if_3_if_and_tmp;
  wire FpAdd_8U_23U_if_3_if_and_tmp_1;
  wire FpAdd_8U_23U_if_3_if_and_tmp_2;
  wire FpAdd_8U_23U_if_3_if_and_tmp_3;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp;
  wire [7:0] z_out_4;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1;
  wire [7:0] z_out_5;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2;
  wire [7:0] z_out_6;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3;
  wire [7:0] z_out_7;
  wire FpAdd_8U_23U_if_2_and_tmp;
  wire [49:0] z_out_12;
  wire FpAdd_8U_23U_if_2_and_tmp_1;
  wire [49:0] z_out_13;
  wire FpAdd_8U_23U_if_2_and_tmp_2;
  wire [49:0] z_out_14;
  wire FpAdd_8U_23U_if_2_and_tmp_3;
  wire [49:0] z_out_15;
  wire chn_alu_in_rsci_ld_core_psct_mx0c0;
  wire alu_loop_op_mux_204_mx1w1;
  wire [21:0] AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0;
  wire [7:0] AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0;
  wire chn_alu_op_rsci_ld_core_psct_mx0c1;
  wire alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
  wire main_stage_v_1_mx0c1;
  wire cfg_alu_src_1_sva_st_1_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0;
  wire alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0;
  wire alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0;
  wire alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0;
  wire alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  wire alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0;
  wire main_stage_v_3_mx0c1;
  wire FpNormalize_8U_49U_if_or_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_1_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_2_itm_mx0w0;
  wire FpNormalize_8U_49U_if_or_3_itm_mx0w0;
  wire main_stage_v_4_mx0c1;
  wire [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0;
  wire [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0;
  wire [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0;
  wire [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0;
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0;
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0;
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0;
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0;
  wire alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1;
  wire FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1;
  wire FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1;
  wire FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1;
  wire alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  wire FpAlu_8U_23U_o_0_sva_2_mx0w0;
  wire AluOut_data_2_0_sva_3_mx0w0;
  wire [31:0] alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0;
  wire [31:0] alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0;
  wire [31:0] alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0;
  wire [31:0] alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0;
  wire alu_loop_op_else_nor_dfs;
  wire FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0;
  wire alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_sva;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_3_sva;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_2_sva;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_1_sva;
  wire FpMantRNE_49U_24U_else_carry_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_3_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_2_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0;
  wire FpMantRNE_49U_24U_else_carry_1_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0;
  wire FpAlu_8U_23U_o_0_lpi_1_dfm_2;
  wire [21:0] FpAlu_8U_23U_o_22_1_lpi_1_dfm_2;
  wire [7:0] FpAlu_8U_23U_o_30_23_lpi_1_dfm_2;
  wire FpAlu_8U_23U_and_30_cse;
  wire FpAlu_8U_23U_and_31_m1c;
  wire FpAlu_8U_23U_and_44_cse;
  wire FpAlu_8U_23U_and_45_cse;
  wire [31:0] alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0;
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_1_sva;
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_1_sva;
  wire [31:0] alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0;
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_2_sva;
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_2_sva;
  wire [31:0] alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0;
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_3_sva;
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_3_sva;
  wire [31:0] alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0;
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_sva;
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_sva;
  wire [30:0] IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1;
  wire [30:0] IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1;
  wire [30:0] IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1;
  wire [30:0] IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1;
  wire [31:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0;
  wire [31:0] FpCmp_8U_23U_false_o_2_lpi_1_dfm_2;
  wire FpAlu_8U_23U_and_48_m1c;
  wire FpAlu_8U_23U_and_52_m1c;
  wire FpAlu_8U_23U_and_56_m1c;
  wire FpAlu_8U_23U_and_40_m1c;
  wire FpNormalize_8U_49U_oelse_not_9;
  wire FpNormalize_8U_49U_oelse_not_11;
  wire FpNormalize_8U_49U_oelse_not_13;
  wire FpNormalize_8U_49U_oelse_not_15;
  wire [7:0] else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23;
  wire [7:0] else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23;
  wire [7:0] else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23;
  wire [30:0] else_AluOp_data_1_lpi_1_dfm_mx2_30_0;
  wire [7:0] else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7;
  wire chn_alu_out_or_cse;
  wire chn_alu_out_and_18_cse;
  wire cfg_alu_algo_cfg_alu_algo_or_3_cse;
  reg reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse;
  wire FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse;
  wire IsNaN_8U_23U_aelse_and_cse;
  wire else_AluOp_data_and_10_cse;
  wire AluIn_data_and_1_cse;
  wire FpAdd_8U_23U_and_39_cse;
  wire FpAdd_8U_23U_int_mant_p1_or_3_cse;
  wire FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse;
  wire nand_109_cse;
  wire nor_430_cse;
  wire and_564_cse;
  wire IsNaN_8U_23U_aelse_and_8_cse;
  wire IsNaN_8U_23U_1_aelse_and_cse;
  wire FpAlu_8U_23U_and_82_cse;
  wire FpCmp_8U_23U_true_o_and_cse;
  wire FpCmp_8U_23U_false_o_and_1_cse;
  wire and_cse;
  wire AluOut_data_and_8_cse;
  wire IntSaturation_33U_32U_and_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_12_cse;
  wire and_550_cse;
  wire IsNaN_8U_23U_aelse_and_12_cse;
  wire FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse;
  wire FpCmp_8U_23U_true_o_and_5_cse;
  wire FpAlu_8U_23U_and_88_cse;
  wire FpCmp_8U_23U_false_o_and_6_cse;
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse;
  wire IntSaturation_33U_32U_and_11_cse;
  wire AluOut_data_and_15_cse;
  wire IsZero_8U_23U_and_6_cse;
  wire IsNaN_8U_23U_aelse_and_16_cse;
  wire AluOut_data_and_17_cse;
  wire FpCmp_8U_23U_true_o_and_9_cse;
  wire FpAlu_8U_23U_and_94_cse;
  wire or_1050_cse;
  wire or_1055_cse;
  wire IntSaturation_33U_32U_if_and_9_cse;
  wire FpAlu_8U_23U_and_102_cse;
  wire AluIn_data_and_cse;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse;
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse;
  wire alu_loop_op_else_else_if_and_cse;
  wire alu_loop_op_else_else_if_and_1_cse;
  reg [1:0] reg_cfg_alu_algo_1_sva_st_13_cse;
  wire FpAdd_8U_23U_is_addition_and_8_cse;
  wire FpAdd_8U_23U_int_mant_p1_and_4_cse;
  wire FpMantRNE_49U_24U_else_and_4_cse;
  wire IsZero_8U_23U_and_4_cse;
  wire AluOut_data_and_12_cse;
  wire FpAlu_8U_23U_or_cse;
  wire IsNaN_8U_23U_2_and_6_cse;
  reg reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse;
  reg reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse;
  reg reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse;
  wire or_dcpl;
  wire mux_tmp;
  wire mux_tmp_348;
  wire mux_tmp_349;
  wire mux_tmp_350;
  wire or_dcpl_272;
  wire FpAdd_8U_23U_and_4_tmp;
  wire FpAdd_8U_23U_and_10_tmp;
  wire FpAdd_8U_23U_and_16_tmp;
  wire FpAdd_8U_23U_and_22_tmp;
  wire nor_437_cse;
  wire and_734_cse;
  wire or_1087_cse;
  wire [1:0] cfg_alu_algo_cfg_alu_algo_mux_3_itm;
  wire alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2;
  wire alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2;
  wire alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2;
  wire alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2;
  wire alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  wire alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1;
  wire alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1;
  wire alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1;
  wire alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1;
  wire alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  wire alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1;
  wire alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1;
  wire alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1;
  wire alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1;
  wire alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1;
  wire FpCmp_8U_23U_true_if_acc_4_itm_8;
  wire FpCmp_8U_23U_true_if_acc_6_itm_8;
  wire FpCmp_8U_23U_false_else_if_acc_6_itm_8;
  wire FpCmp_8U_23U_true_else_else_if_acc_4_itm_23;
  wire FpCmp_8U_23U_true_if_acc_8_itm_8;
  wire FpCmp_8U_23U_true_if_acc_10_itm_8;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1;
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1;
  wire mux_281_cse;
  wire IsNaN_8U_23U_2_and_9_cse;

  wire[0:0] oWidth_iWidth_prb;
  wire[0:0] oWidth_iWidth_prb_1;
  wire[0:0] oWidth_iWidth_prb_2;
  wire[0:0] oWidth_iWidth_prb_3;
  wire[0:0] alu_loop_op_mux_209_nl;
  wire[0:0] FpAlu_8U_23U_mux1h_147_nl;
  wire[21:0] FpAlu_8U_23U_and_5_nl;
  wire[21:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_nl;
  wire[0:0] FpAlu_8U_23U_not_24_nl;
  wire[7:0] FpAlu_8U_23U_and_4_nl;
  wire[7:0] FpAlu_8U_23U_mux1h_145_nl;
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_nl;
  wire[0:0] FpAdd_8U_23U_and_6_nl;
  wire[0:0] FpAdd_8U_23U_and_28_nl;
  wire[0:0] FpAdd_8U_23U_and_9_nl;
  wire[0:0] FpAlu_8U_23U_not_27_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] alu_loop_op_mux_210_nl;
  wire[0:0] FpAlu_8U_23U_mux1h_151_nl;
  wire[21:0] FpAlu_8U_23U_and_8_nl;
  wire[21:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl;
  wire[0:0] FpAlu_8U_23U_not_23_nl;
  wire[7:0] FpAlu_8U_23U_and_7_nl;
  wire[7:0] FpAlu_8U_23U_mux1h_149_nl;
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl;
  wire[0:0] FpAdd_8U_23U_and_29_nl;
  wire[0:0] FpAdd_8U_23U_and_13_nl;
  wire[0:0] FpAdd_8U_23U_and_30_nl;
  wire[0:0] FpAdd_8U_23U_and_15_nl;
  wire[0:0] FpAlu_8U_23U_not_26_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] alu_loop_op_mux_212_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] nand_nl;
  wire[0:0] and_502_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] nand_18_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] or_43_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] else_AluOp_data_else_AluOp_data_nor_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] nor_350_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] and_500_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] nor_339_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] and_499_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] nor_332_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] nor_314_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] and_498_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] nor_317_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] nor_319_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_320_nl;
  wire[0:0] nor_322_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] and_497_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] nor_310_nl;
  wire[0:0] nor_311_nl;
  wire[0:0] nor_312_nl;
  wire[0:0] nor_313_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] or_182_nl;
  wire[0:0] or_962_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] nor_309_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] nor_302_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] nor_300_nl;
  wire[22:0] else_AluOp_data_else_AluOp_data_mux_7_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl;
  wire[22:0] alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl;
  wire[23:0] nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl;
  wire[0:0] FpAdd_8U_23U_is_inf_mux_3_nl;
  wire[0:0] and_192_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] nor_290_nl;
  wire[0:0] nor_291_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] nor_293_nl;
  wire[0:0] or_225_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] or_239_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] or_236_nl;
  wire[22:0] else_AluOp_data_else_AluOp_data_mux_6_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl;
  wire[22:0] alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[23:0] nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl;
  wire[0:0] FpAdd_8U_23U_is_inf_mux_2_nl;
  wire[0:0] and_196_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] or_741_nl;
  wire[0:0] mux_329_nl;
  wire[22:0] else_AluOp_data_else_AluOp_data_mux_5_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl;
  wire[22:0] alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl;
  wire[23:0] nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl;
  wire[0:0] FpAdd_8U_23U_is_inf_mux_1_nl;
  wire[0:0] and_200_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] or_744_nl;
  wire[0:0] mux_331_nl;
  wire[22:0] else_AluOp_data_else_AluOp_data_mux_4_nl;
  wire[22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl;
  wire[22:0] alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  wire[0:0] FpAdd_8U_23U_is_inf_mux_nl;
  wire[0:0] and_204_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] or_747_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] or_270_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] or_273_nl;
  wire[0:0] or_275_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] or_1100_nl;
  wire[0:0] or_1106_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] or_280_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] or_288_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] nor_272_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] nor_270_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] or_299_nl;
  wire[0:0] or_301_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] or_304_nl;
  wire[0:0] or_307_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] or_312_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] nor_267_nl;
  wire[0:0] nor_268_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] and_218_nl;
  wire[0:0] and_220_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] or_1046_nl;
  wire[0:0] mux_nl;
  wire[0:0] or_1048_nl;
  wire[0:0] and_729_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] or_333_nl;
  wire[0:0] and_496_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] or_334_nl;
  wire[0:0] and_495_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] or_335_nl;
  wire[0:0] and_494_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] or_336_nl;
  wire[0:0] and_493_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] nor_263_nl;
  wire[0:0] nor_265_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] nor_260_nl;
  wire[0:0] nor_262_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] nor_259_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] nor_254_nl;
  wire[0:0] nor_256_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] or_961_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] nor_251_nl;
  wire[0:0] or_960_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] or_959_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] or_958_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] nand_29_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] or_400_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] nor_241_nl;
  wire[0:0] nor_243_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_or_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] or_422_nl;
  wire[0:0] or_420_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] or_426_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_or_3_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_or_2_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_or_1_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] or_438_nl;
  wire[0:0] or_440_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] or_441_nl;
  wire[0:0] or_443_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] or_446_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] or_444_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] or_450_nl;
  wire[0:0] nor_80_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] or_453_nl;
  wire[0:0] nor_81_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] nor_237_nl;
  wire[0:0] nor_238_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] or_463_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] nor_232_nl;
  wire[0:0] nor_233_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] nor_227_nl;
  wire[0:0] nor_228_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] nor_222_nl;
  wire[0:0] nor_223_nl;
  wire[0:0] FpAlu_8U_23U_and_9_nl;
  wire[0:0] FpAlu_8U_23U_and_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] nor_219_nl;
  wire[0:0] nor_220_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] nor_217_nl;
  wire[0:0] nor_218_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] nor_215_nl;
  wire[0:0] nor_216_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] nor_213_nl;
  wire[0:0] nor_214_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] and_485_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] nor_208_nl;
  wire[0:0] nor_210_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] nor_207_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] nor_206_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] and_478_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] nor_204_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] nor_205_nl;
  wire[0:0] AluOut_data_or_1_nl;
  wire[0:0] alu_loop_op_else_mux_1_nl;
  wire[0:0] AluOut_data_or_2_nl;
  wire[0:0] alu_loop_op_else_mux_2_nl;
  wire[0:0] AluOut_data_and_7_nl;
  wire[0:0] alu_loop_op_else_mux_nl;
  wire[0:0] AluOut_data_or_nl;
  wire[0:0] FpAlu_8U_23U_mux_21_nl;
  wire[0:0] AluOut_data_or_3_nl;
  wire[0:0] FpAlu_8U_23U_mux_20_nl;
  wire[0:0] AluOut_data_and_3_nl;
  wire[0:0] alu_loop_op_else_mux_3_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] nor_203_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] nor_200_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] nor_195_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] nor_192_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] or_1069_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] or_1076_nl;
  wire[0:0] FpAlu_8U_23U_mux1h_144_nl;
  wire[0:0] FpAlu_8U_23U_or_145_nl;
  wire[0:0] FpAlu_8U_23U_or_146_nl;
  wire[0:0] FpAlu_8U_23U_mux1h_148_nl;
  wire[0:0] FpAlu_8U_23U_or_147_nl;
  wire[0:0] FpAlu_8U_23U_or_148_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] FpAlu_8U_23U_and_74_nl;
  wire[0:0] FpAlu_8U_23U_and_75_nl;
  wire[0:0] FpAlu_8U_23U_and_76_nl;
  wire[0:0] FpAlu_8U_23U_and_77_nl;
  wire[0:0] FpAlu_8U_23U_and_80_nl;
  wire[0:0] alu_loop_op_else_mux_5_nl;
  wire[0:0] FpAlu_8U_23U_and_81_nl;
  wire[0:0] alu_loop_op_else_mux_4_nl;
  wire[0:0] FpAlu_8U_23U_and_66_nl;
  wire[0:0] FpAlu_8U_23U_and_67_nl;
  wire[0:0] FpAlu_8U_23U_and_68_nl;
  wire[0:0] FpAlu_8U_23U_and_69_nl;
  wire[0:0] FpAlu_8U_23U_and_72_nl;
  wire[0:0] FpAlu_8U_23U_and_73_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] and_74_nl;
  wire[0:0] nand_30_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] or_624_nl;
  wire[0:0] or_619_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] nand_35_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nor_178_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] nor_176_nl;
  wire[0:0] nand_38_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] FpAlu_8U_23U_mux1h_155_nl;
  wire[21:0] FpAlu_8U_23U_and_11_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_154_nl;
  wire[0:0] FpAlu_8U_23U_not_22_nl;
  wire[7:0] FpAlu_8U_23U_and_10_nl;
  wire[7:0] FpAlu_8U_23U_mux1h_153_nl;
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl;
  wire[0:0] FpAdd_8U_23U_and_31_nl;
  wire[0:0] FpAdd_8U_23U_and_19_nl;
  wire[0:0] FpAdd_8U_23U_and_32_nl;
  wire[0:0] FpAdd_8U_23U_and_21_nl;
  wire[0:0] FpAlu_8U_23U_not_25_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] and_97_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_38_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_39_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_40_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_41_nl;
  wire[8:0] acc_nl;
  wire[9:0] nl_acc_nl;
  wire[5:0] FpNormalize_8U_49U_else_mux_4_nl;
  wire[0:0] nor_436_nl;
  wire[8:0] acc_1_nl;
  wire[9:0] nl_acc_1_nl;
  wire[5:0] FpNormalize_8U_49U_else_mux_5_nl;
  wire[0:0] nor_435_nl;
  wire[8:0] acc_2_nl;
  wire[9:0] nl_acc_2_nl;
  wire[5:0] FpNormalize_8U_49U_else_mux_6_nl;
  wire[0:0] nor_434_nl;
  wire[8:0] acc_3_nl;
  wire[9:0] nl_acc_3_nl;
  wire[5:0] FpNormalize_8U_49U_else_mux_7_nl;
  wire[0:0] nor_433_nl;
  wire[31:0] alu_loop_op_else_alu_loop_op_else_mux_3_nl;
  wire[0:0] alu_loop_op_else_not_18_nl;
  wire[31:0] alu_loop_op_else_alu_loop_op_else_mux_2_nl;
  wire[0:0] alu_loop_op_else_not_20_nl;
  wire[2:0] alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl;
  wire[3:0] nl_alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl;
  wire[31:0] alu_loop_op_else_alu_loop_op_else_mux_1_nl;
  wire[0:0] alu_loop_op_else_not_22_nl;
  wire[31:0] alu_loop_op_else_alu_loop_op_else_mux_nl;
  wire[0:0] alu_loop_op_else_not_21_nl;
  wire[2:0] alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl;
  wire[3:0] nl_alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl;
  wire[2:0] alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl;
  wire[3:0] nl_alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl;
  wire[2:0] alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl;
  wire[3:0] nl_alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl;
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl;
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl;
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  wire[21:0] FpAlu_8U_23U_mux1h_35_nl;
  wire[0:0] FpAlu_8U_23U_not_21_nl;
  wire[7:0] FpAlu_8U_23U_mux1h_34_nl;
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl;
  wire[0:0] FpAdd_8U_23U_and_33_nl;
  wire[0:0] FpAdd_8U_23U_and_25_nl;
  wire[0:0] FpAdd_8U_23U_and_34_nl;
  wire[0:0] FpAdd_8U_23U_and_27_nl;
  wire[0:0] FpAlu_8U_23U_and_62_nl;
  wire[0:0] FpAlu_8U_23U_not_17_nl;
  wire[33:0] acc_8_nl;
  wire[34:0] nl_acc_8_nl;
  wire[31:0] alu_loop_op_else_if_mux_8_nl;
  wire[31:0] alu_loop_op_else_if_mux_9_nl;
  wire[33:0] acc_10_nl;
  wire[34:0] nl_acc_10_nl;
  wire[31:0] alu_loop_op_else_if_mux_12_nl;
  wire[31:0] alu_loop_op_else_if_mux_13_nl;
  wire[33:0] acc_11_nl;
  wire[34:0] nl_acc_11_nl;
  wire[31:0] alu_loop_op_else_if_mux_14_nl;
  wire[31:0] alu_loop_op_else_if_mux_15_nl;
  wire[33:0] acc_9_nl;
  wire[34:0] nl_acc_9_nl;
  wire[31:0] alu_loop_op_else_if_mux_10_nl;
  wire[31:0] alu_loop_op_else_if_mux_11_nl;
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl;
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl;
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl;
  wire[0:0] IntSaturation_33U_32U_and_3_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl;
  wire[0:0] IntSaturation_33U_32U_and_7_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl;
  wire[0:0] IntSaturation_33U_32U_and_5_nl;
  wire[0:0] IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl;
  wire[0:0] IntSaturation_33U_32U_and_1_nl;
  wire[2:0] alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl;
  wire[3:0] nl_alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl;
  wire[2:0] alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl;
  wire[3:0] nl_alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl;
  wire[2:0] alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl;
  wire[3:0] nl_alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl;
  wire[2:0] alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl;
  wire[3:0] nl_alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_4_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_4_nl;
  wire[23:0] FpCmp_8U_23U_true_else_else_if_acc_8_nl;
  wire[25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_8_nl;
  wire[0:0] asn_FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_nor_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] nor_168_nl;
  wire[0:0] and_446_nl;
  wire[0:0] asn_FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_nor_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] or_864_nl;
  wire[23:0] FpCmp_8U_23U_true_else_else_if_acc_7_nl;
  wire[25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_7_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_8_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_8_nl;
  wire[0:0] asn_FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_nor_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] nor_165_nl;
  wire[0:0] and_444_nl;
  wire[23:0] FpCmp_8U_23U_true_else_else_if_acc_6_nl;
  wire[25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_6_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_10_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_10_nl;
  wire[0:0] asn_FpCmp_8U_23U_true_o_lpi_1_dfm_1_nor_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] nor_163_nl;
  wire[0:0] and_443_nl;
  wire[0:0] or_876_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] and_336_nl;
  wire[0:0] nor_162_nl;
  wire[0:0] or_880_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] and_338_nl;
  wire[0:0] nor_159_nl;
  wire[0:0] or_884_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] and_340_nl;
  wire[0:0] nor_156_nl;
  wire[0:0] FpAlu_8U_23U_and_61_nl;
  wire[0:0] FpCmp_8U_23U_false_mux_4_nl;
  wire[0:0] FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_nl;
  wire[0:0] FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_nl;
  wire[8:0] alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  wire[8:0] alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl;
  wire[10:0] nl_alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl;
  wire[8:0] alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl;
  wire[10:0] nl_alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl;
  wire[8:0] alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl;
  wire[10:0] nl_alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_4_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_4_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_6_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_6_nl;
  wire[8:0] FpCmp_8U_23U_false_else_if_acc_6_nl;
  wire[10:0] nl_FpCmp_8U_23U_false_else_if_acc_6_nl;
  wire[23:0] FpCmp_8U_23U_true_else_else_if_acc_4_nl;
  wire[25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_4_nl;
  wire[22:0] else_else_mux_13_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_8_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_8_nl;
  wire[8:0] FpCmp_8U_23U_true_if_acc_10_nl;
  wire[10:0] nl_FpCmp_8U_23U_true_if_acc_10_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] or_967_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] or_965_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] nor_357_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] or_87_nl;
  wire[0:0] or_230_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] or_233_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] or_323_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] or_386_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] or_383_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] or_417_nl;
  wire[0:0] or_419_nl;
  wire[0:0] or_428_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] or_432_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_474_nl;
  wire[0:0] nor_187_nl;
  wire[0:0] or_609_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] or_601_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] or_607_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] or_610_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] or_612_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] or_629_nl;
  wire[0:0] nor_117_nl;
  wire[0:0] nor_124_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] nor_143_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  wire[8:0] acc_4_nl;
  wire[9:0] nl_acc_4_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_15_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_16_nl;
  wire[8:0] acc_5_nl;
  wire[9:0] nl_acc_5_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_17_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_18_nl;
  wire[8:0] acc_6_nl;
  wire[9:0] nl_acc_6_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_19_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_20_nl;
  wire[8:0] acc_7_nl;
  wire[9:0] nl_acc_7_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_21_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_22_nl;
  wire[50:0] acc_12_nl;
  wire[51:0] nl_acc_12_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_8_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_9_nl;
  wire[50:0] acc_13_nl;
  wire[51:0] nl_acc_13_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_10_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_11_nl;
  wire[50:0] acc_14_nl;
  wire[51:0] nl_acc_14_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_12_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_13_nl;
  wire[50:0] acc_15_nl;
  wire[51:0] nl_acc_15_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_14_nl;
  wire[48:0] FpAdd_8U_23U_else_2_mux_15_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2
      , (else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0])};
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl = nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl[7:0];
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {(alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_a;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_a = {alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2
      , (else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0])};
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl;
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl = nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl[7:0];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s = {(alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = {alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2
      , (else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0])};
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl;
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl = nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl[7:0];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s = {(alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_a;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_a = {alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2
      , (else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0])};
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl;
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl = nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl[7:0];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s = {(alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_a;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_a = {alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_128[118:96])};
  wire[7:0] alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl;
  wire[8:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl;
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl = nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl[7:0];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s = {(alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = {alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5
      , (AluIn_data_sva_128[86:64])};
  wire[7:0] alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl;
  wire[8:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl;
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl = nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl[7:0];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s = {(alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_a;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_a = {alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4
      , (AluIn_data_sva_128[54:32])};
  wire[7:0] alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl;
  wire[8:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl;
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl = nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl[7:0];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s = {(alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5[0]))};
  wire [23:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3
      , (AluIn_data_sva_128[22:0])};
  wire[7:0] alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire[8:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5[7:1]))})
      + 8'b1101;
  assign alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl = nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl[7:0];
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {(alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5[0]))};
  wire [48:0] nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa;
  assign nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_2_leading_sign_49_0_2_rg_mantissa;
  assign nl_alu_loop_op_2_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_3_leading_sign_49_0_1_rg_mantissa;
  assign nl_alu_loop_op_3_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_4_leading_sign_49_0_3_rg_mantissa;
  assign nl_alu_loop_op_4_leading_sign_49_0_3_rg_mantissa = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg_a;
  assign nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg_a = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg_a;
  assign nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg_a;
  assign nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg_a = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0];
  wire [48:0] nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0];
  wire [127:0] nl_Y_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d;
  assign nl_Y_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d = {chn_alu_out_rsci_d_127
      , chn_alu_out_rsci_d_126_119 , chn_alu_out_rsci_d_118_97 , chn_alu_out_rsci_d_96
      , chn_alu_out_rsci_d_95 , chn_alu_out_rsci_d_94_87 , chn_alu_out_rsci_d_86_65
      , chn_alu_out_rsci_d_64 , chn_alu_out_rsci_d_63 , chn_alu_out_rsci_d_62_55
      , chn_alu_out_rsci_d_54_33 , chn_alu_out_rsci_d_32 , chn_alu_out_rsci_d_31
      , chn_alu_out_rsci_d_30_23 , chn_alu_out_rsci_d_22_1 , chn_alu_out_rsci_d_0};
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_19_mx0w1)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg (
      .a(nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_a[23:0]),
      .s(nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_13_mx0w1)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_7_mx0w1)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg (
      .a(nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_a[23:0]),
      .s(nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_1_mx0w1)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg (
      .a(nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_a[23:0]),
      .s(nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_sva)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
      .a(nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a[23:0]),
      .s(nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_3_sva)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg (
      .a(nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_a[23:0]),
      .s(nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_2_sva)
    );
  SDP_Y_CORE_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_1_sva)
    );
  SDP_Y_CORE_leading_sign_49_0  alu_loop_op_1_leading_sign_49_0_rg (
      .mantissa(nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4)
    );
  SDP_Y_CORE_leading_sign_49_0  alu_loop_op_2_leading_sign_49_0_2_rg (
      .mantissa(nl_alu_loop_op_2_leading_sign_49_0_2_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5)
    );
  SDP_Y_CORE_leading_sign_49_0  alu_loop_op_3_leading_sign_49_0_1_rg (
      .mantissa(nl_alu_loop_op_3_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6)
    );
  SDP_Y_CORE_leading_sign_49_0  alu_loop_op_4_leading_sign_49_0_3_rg (
      .mantissa(nl_alu_loop_op_4_leading_sign_49_0_3_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7)
    );
  SDP_Y_CORE_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg (
      .a(nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7),
      .z(alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_itm)
    );
  SDP_Y_CORE_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg (
      .a(nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6),
      .z(alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_itm)
    );
  SDP_Y_CORE_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg (
      .a(nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5),
      .z(alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_itm)
    );
  SDP_Y_CORE_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4),
      .z(alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci Y_alu_core_chn_alu_in_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsc_z(chn_alu_in_rsc_z),
      .chn_alu_in_rsc_vz(chn_alu_in_rsc_vz),
      .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_alu_in_rsci_iswt0(chn_alu_in_rsci_iswt0),
      .chn_alu_in_rsci_bawt(chn_alu_in_rsci_bawt),
      .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
      .chn_alu_in_rsci_ld_core_psct(chn_alu_in_rsci_ld_core_psct),
      .chn_alu_in_rsci_d_mxwt(chn_alu_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci Y_alu_core_chn_alu_op_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
      .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
      .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_op_rsci_iswt0(chn_alu_op_rsci_iswt0),
      .chn_alu_op_rsci_bawt(chn_alu_op_rsci_bawt),
      .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
      .chn_alu_op_rsci_ld_core_psct(chn_alu_op_rsci_ld_core_psct),
      .chn_alu_op_rsci_d_mxwt(chn_alu_op_rsci_d_mxwt)
    );
  SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci Y_alu_core_chn_alu_out_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_out_rsc_z(chn_alu_out_rsc_z),
      .chn_alu_out_rsc_vz(chn_alu_out_rsc_vz),
      .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_alu_out_rsci_iswt0(chn_alu_out_rsci_iswt0),
      .chn_alu_out_rsci_bawt(chn_alu_out_rsci_bawt),
      .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp),
      .chn_alu_out_rsci_ld_core_psct(reg_chn_alu_out_rsci_ld_core_psct_cse),
      .chn_alu_out_rsci_d(nl_Y_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d[127:0])
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz),
      .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_bypass_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_bypass_rsc_triosy_obj_bawt(cfg_alu_bypass_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj Y_alu_core_cfg_alu_src_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz),
      .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_src_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_src_rsc_triosy_obj_bawt(cfg_alu_src_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj Y_alu_core_cfg_alu_op_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz),
      .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_op_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_op_rsc_triosy_obj_bawt(cfg_alu_op_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj Y_alu_core_cfg_alu_algo_rsc_triosy_obj_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz),
      .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .cfg_alu_algo_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
      .cfg_alu_algo_rsc_triosy_obj_bawt(cfg_alu_algo_rsc_triosy_obj_bawt)
    );
  SDP_Y_CORE_Y_alu_core_staller Y_alu_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
      .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp)
    );
  SDP_Y_CORE_Y_alu_core_core_fsm Y_alu_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign oWidth_iWidth_prb = alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
  // assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
  // PSL alu_loop_op_1_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_1 = alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
  // assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
  // PSL alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1 : assert { oWidth_iWidth_prb_1 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_2 = alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
  // assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
  // PSL alu_loop_op_3_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb_2 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_3 = alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
  // assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
  // PSL alu_loop_op_4_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1 : assert { oWidth_iWidth_prb_3 } @rose(nvdla_core_clk);
  assign chn_alu_out_or_cse = (and_dcpl_37 & or_1087_cse) | and_dcpl_40;
  assign chn_alu_out_and_cse = core_wen & chn_alu_out_or_cse;
  assign chn_alu_out_and_1_cse = core_wen & (~ or_dcpl_23);
  assign nor_437_cse = ~(asn_267 | or_dcpl);
  assign or_1087_cse = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt;
  assign and_734_cse = (or_dcpl_272 | FpAlu_8U_23U_nor_dfs_6 | FpAlu_8U_23U_equal_tmp_23
      | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8) & or_1087_cse
      & main_stage_v_4 & core_wen;
  assign chn_alu_out_and_8_cse = core_wen & (~ (fsm_output[0]));
  assign chn_alu_out_and_18_cse = chn_alu_out_and_8_cse & (~ or_dcpl_23);
  assign nand_nl = ~(or_937_cse & (~(nor_269_cse | chn_alu_in_rsci_bawt | (~ and_dcpl_4))));
  assign and_502_nl = or_1087_cse & chn_alu_in_rsci_bawt;
  assign mux_15_nl = MUX_s_1_2_2((and_502_nl), (nand_nl), main_stage_v_1);
  assign AluIn_data_and_cse = core_wen & (~ or_dcpl_49) & (mux_15_nl);
  assign nor_6_cse = ~((cfg_precision!=2'b10));
  assign nor_5_cse = ~(cfg_alu_bypass_rsci_d | (~ chn_alu_in_rsci_bawt));
  assign or_28_cse = (cfg_alu_algo_1_sva_st_20!=2'b01) | (cfg_alu_algo_1_sva_st[1]);
  assign cfg_alu_algo_cfg_alu_algo_or_3_cse = (or_dcpl_14 & and_dcpl_78) | and_dcpl_81;
  assign cfg_alu_algo_cfg_alu_algo_mux_3_itm = MUX_v_2_2_2(cfg_alu_algo_rsci_d, cfg_alu_algo_1_sva_st_20,
      and_dcpl_81);
  assign or_937_cse = (~ cfg_alu_src_1_sva_st_1) | chn_alu_op_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign or_963_cse = (~ cfg_alu_src_1_sva_st_1) | chn_alu_op_rsci_bawt;
  assign and_501_cse = or_963_cse & cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_167_rgt = or_tmp_386 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1
      & alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign IsNaN_8U_23U_aelse_and_cse = core_wen & (~ and_dcpl_32) & not_tmp_29;
  assign FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse = and_dcpl_78
      | and_dcpl_99;
  assign FpAdd_8U_23U_is_addition_and_8_cse = core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
      & not_tmp_29;
  assign nor_367_nl = ~((~ main_stage_v_1) | io_read_cfg_alu_bypass_rsc_svs_st_1
      | (~(cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt &
      cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt & or_963_cse)));
  assign nor_368_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5);
  assign mux_43_nl = MUX_s_1_2_2((nor_368_nl), (nor_367_nl), or_1087_cse);
  assign else_AluOp_data_and_10_cse = core_wen & (~ and_dcpl_32) & (mux_43_nl);
  assign mux_44_nl = MUX_s_1_2_2(main_stage_v_2, and_dcpl_4, or_1087_cse);
  assign mux_45_nl = MUX_s_1_2_2(not_tmp_38, (mux_44_nl), or_937_cse);
  assign mux_46_nl = MUX_s_1_2_2(not_tmp_38, (mux_45_nl), main_stage_v_1);
  assign AluIn_data_and_1_cse = core_wen & (~ and_dcpl_32) & (mux_46_nl);
  assign FpAdd_8U_23U_and_39_cse = core_wen & (~ and_dcpl_32) & not_tmp_57;
  assign FpAdd_8U_23U_int_mant_p1_or_3_cse = or_dcpl_86 | and_dcpl_99;
  assign FpAdd_8U_23U_int_mant_p1_and_4_cse = core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
      & not_tmp_57;
  assign and_550_cse = core_wen & (~ and_dcpl_32) & mux_tmp_53;
  assign nor_33_cse = ~(alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49])));
  assign FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse = (or_1087_cse & (~ alu_loop_op_unequal_tmp_7))
      | and_dcpl_108;
  assign nor_37_cse = ~(alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1 | (~ (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49])));
  assign nor_41_cse = ~(alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1 | (~ (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49])));
  assign nor_45_cse = ~(alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1 | (~ (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49])));
  assign nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_sva);
  assign alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl = nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl[22:0];
  assign FpAdd_8U_23U_is_inf_mux_3_nl = MUX_s_1_2_2(nor_45_cse, FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0,
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp);
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl = MUX_v_23_2_2((alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl),
      23'b11111111111111111111111, (FpAdd_8U_23U_is_inf_mux_3_nl));
  assign and_192_nl = or_1087_cse & (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8);
  assign else_AluOp_data_else_AluOp_data_mux_7_nl = MUX_v_23_2_2(else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2,
      (FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl), and_192_nl);
  assign or_735_nl = IsNaN_8U_23U_land_lpi_1_dfm_11 | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_8;
  assign mux_327_nl = MUX_s_1_2_2(mux_tmp_311, or_tmp_657, IsNaN_8U_23U_land_lpi_1_dfm_11);
  assign mux_328_nl = MUX_s_1_2_2((mux_327_nl), (or_735_nl), IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign AluIn_data_mux1h_7_itm = MUX_v_31_2_2(({8'b0 , (else_AluOp_data_else_AluOp_data_mux_7_nl)}),
      AluIn_data_sva_3_126_96_1, mux_328_nl);
  assign nand_109_cse = ~((~((cfg_alu_algo_1_sva_st_24==2'b10))) & FpAlu_8U_23U_equal_tmp_22);
  assign nor_430_cse = ~(alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_st_6);
  assign and_564_cse = (cfg_alu_algo_1_sva_st_24==2'b10);
  assign nor_290_nl = ~((cfg_alu_algo_1_sva_st_24!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_5)
      | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | io_read_cfg_alu_bypass_rsc_svs_7
      | alu_loop_op_unequal_tmp_7);
  assign nor_291_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7);
  assign mux_105_nl = MUX_s_1_2_2((nor_291_nl), (nor_290_nl), FpAlu_8U_23U_equal_tmp_22);
  assign nor_293_nl = ~((cfg_alu_algo_1_sva_st_25[1]) | (~ FpAlu_8U_23U_equal_tmp_23));
  assign or_225_nl = (~ FpAlu_8U_23U_nor_dfs_6) | (cfg_alu_algo_1_sva_st_25[0]);
  assign mux_106_nl = MUX_s_1_2_2((nor_293_nl), FpAlu_8U_23U_equal_tmp_23, or_225_nl);
  assign nor_292_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8
      | io_read_cfg_alu_bypass_rsc_svs_st_7 | (mux_106_nl));
  assign mux_107_nl = MUX_s_1_2_2((nor_292_nl), (mux_105_nl), or_1087_cse);
  assign IsNaN_8U_23U_aelse_and_8_cse = core_wen & (~ and_dcpl_32) & (mux_107_nl);
  assign IsNaN_8U_23U_1_aelse_and_cse = core_wen & (~ and_dcpl_32) & (~ mux_109_itm);
  assign or_239_nl = nor_269_cse | (cfg_alu_algo_1_sva_st_24!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_110_nl = MUX_s_1_2_2(or_tmp_224, or_tmp_75, or_1087_cse);
  assign or_236_nl = (cfg_alu_algo_1_sva_st_25!=2'b10);
  assign mux_111_nl = MUX_s_1_2_2((mux_110_nl), (or_239_nl), or_236_nl);
  assign FpMantRNE_49U_24U_else_and_4_cse = core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
      & (~ (mux_111_nl));
  assign nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_3_sva);
  assign alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl = nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl[22:0];
  assign FpAdd_8U_23U_is_inf_mux_2_nl = MUX_s_1_2_2(nor_41_cse, FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0,
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp);
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl = MUX_v_23_2_2((alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl),
      23'b11111111111111111111111, (FpAdd_8U_23U_is_inf_mux_2_nl));
  assign and_196_nl = or_1087_cse & (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8);
  assign else_AluOp_data_else_AluOp_data_mux_6_nl = MUX_v_23_2_2(else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2,
      (FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl), and_196_nl);
  assign or_741_nl = IsNaN_8U_23U_land_3_lpi_1_dfm_11 | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_8;
  assign mux_329_nl = MUX_s_1_2_2(mux_tmp_311, or_tmp_657, IsNaN_8U_23U_land_3_lpi_1_dfm_11);
  assign mux_330_nl = MUX_s_1_2_2((mux_329_nl), (or_741_nl), IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign AluIn_data_mux1h_9_itm = MUX_v_31_2_2(({8'b0 , (else_AluOp_data_else_AluOp_data_mux_6_nl)}),
      AluIn_data_sva_3_94_64_1, mux_330_nl);
  assign nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_2_sva);
  assign alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl = nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl[22:0];
  assign FpAdd_8U_23U_is_inf_mux_1_nl = MUX_s_1_2_2(nor_37_cse, FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0,
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp);
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl = MUX_v_23_2_2((alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl),
      23'b11111111111111111111111, (FpAdd_8U_23U_is_inf_mux_1_nl));
  assign and_200_nl = or_1087_cse & (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8);
  assign else_AluOp_data_else_AluOp_data_mux_5_nl = MUX_v_23_2_2(else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2,
      (FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl), and_200_nl);
  assign or_744_nl = IsNaN_8U_23U_land_2_lpi_1_dfm_11 | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_8;
  assign mux_331_nl = MUX_s_1_2_2(mux_tmp_311, or_tmp_657, IsNaN_8U_23U_land_2_lpi_1_dfm_11);
  assign mux_332_nl = MUX_s_1_2_2((mux_331_nl), (or_744_nl), IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign AluIn_data_mux1h_11_itm = MUX_v_31_2_2(({8'b0 , (else_AluOp_data_else_AluOp_data_mux_5_nl)}),
      AluIn_data_sva_3_62_32_1, mux_332_nl);
  assign nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_1_sva);
  assign alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl = nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_is_inf_mux_nl = MUX_s_1_2_2(nor_33_cse, FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0,
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp);
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl = MUX_v_23_2_2((alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, (FpAdd_8U_23U_is_inf_mux_nl));
  assign and_204_nl = or_1087_cse & (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8);
  assign else_AluOp_data_else_AluOp_data_mux_4_nl = MUX_v_23_2_2(else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2,
      (FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl), and_204_nl);
  assign or_747_nl = IsNaN_8U_23U_land_1_lpi_1_dfm_11 | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_8;
  assign mux_333_nl = MUX_s_1_2_2(mux_tmp_311, or_tmp_657, IsNaN_8U_23U_land_1_lpi_1_dfm_11);
  assign mux_334_nl = MUX_s_1_2_2((mux_333_nl), (or_747_nl), IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign AluIn_data_mux1h_13_itm = MUX_v_31_2_2(({8'b0 , (else_AluOp_data_else_AluOp_data_mux_4_nl)}),
      AluIn_data_sva_3_30_0_1, mux_334_nl);
  assign or_270_nl = alu_loop_op_unequal_tmp_8 | io_read_cfg_alu_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_124_nl = MUX_s_1_2_2((or_270_nl), or_tmp_251, or_1087_cse);
  assign FpAlu_8U_23U_and_82_cse = core_wen & (~ and_dcpl_32) & (~ (mux_124_nl));
  assign or_273_nl = (~ FpAlu_8U_23U_equal_tmp_26) | alu_loop_op_unequal_tmp_8 |
      io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_125_nl = MUX_s_1_2_2((or_273_nl), or_tmp_251, or_1087_cse);
  assign or_275_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ FpAlu_8U_23U_equal_tmp_26) | alu_loop_op_unequal_tmp_8 | io_read_cfg_alu_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign mux_126_nl = MUX_s_1_2_2((or_275_nl), (mux_125_nl), FpAlu_8U_23U_equal_tmp_25);
  assign FpCmp_8U_23U_true_o_and_cse = core_wen & (~ and_dcpl_32) & (~ (mux_126_nl));
  assign and_211_rgt = or_1087_cse & (~ alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp);
  assign or_288_nl = (~ FpAlu_8U_23U_equal_tmp_29) | alu_loop_op_unequal_tmp_8 |
      io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_129_nl = MUX_s_1_2_2((or_288_nl), or_tmp_269, or_1087_cse);
  assign FpCmp_8U_23U_false_o_and_1_cse = core_wen & (~ and_dcpl_32) & (~ (mux_129_nl));
  assign and_213_rgt = or_1087_cse & (~ alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp);
  assign and_215_rgt = or_1087_cse & (~ alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp);
  assign nor_269_cse = ~((~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt);
  assign nor_397_cse = ~(alu_loop_op_unequal_tmp_8 | io_read_cfg_alu_bypass_rsc_svs_8);
  assign and_524_cse = (FpAlu_8U_23U_equal_tmp_29 | FpAlu_8U_23U_equal_tmp_26 | FpAlu_8U_23U_nor_dfs_6
      | FpAlu_8U_23U_equal_tmp_23) & or_1087_cse & nor_397_cse & main_stage_v_4 &
      core_wen;
  assign and_217_rgt = or_1087_cse & (~ alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp);
  assign mux_140_nl = MUX_s_1_2_2(main_stage_v_4, main_stage_v_3, or_1087_cse);
  assign and_cse = core_wen & (~ and_dcpl_32) & (mux_140_nl);
  assign AluOut_data_and_8_cse = core_wen & (~ and_dcpl_32) & (~ mux_143_itm);
  assign mux_144_nl = MUX_s_1_2_2(or_tmp_309, or_tmp_312, or_1087_cse);
  assign IntSaturation_33U_32U_and_cse = core_wen & (~ and_dcpl_32) & (~ (mux_144_nl));
  assign FpMantRNE_49U_24U_else_and_cse = core_wen & (~ or_dcpl_85);
  assign nor_264_cse = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6);
  assign FpAdd_8U_23U_int_mant_p1_and_cse = core_wen & (~(or_dcpl_91 | and_dcpl_32
      | io_read_cfg_alu_bypass_rsc_svs_st_5));
  assign FpAdd_8U_23U_int_mant_p1_and_12_cse = FpAdd_8U_23U_int_mant_p1_and_cse &
      (~ or_dcpl_86);
  assign FpAdd_8U_23U_if_3_and_cse = core_wen & (~ or_dcpl_89);
  assign mux_164_nl = MUX_s_1_2_2(not_tmp_157, nand_tmp_13, or_381_cse);
  assign mux_165_nl = MUX_s_1_2_2(not_tmp_157, nand_tmp_13, or_391_cse);
  assign mux_166_nl = MUX_s_1_2_2((mux_165_nl), (mux_164_nl), nor_6_cse);
  assign mux_167_nl = MUX_s_1_2_2(nand_tmp_13, (mux_166_nl), nor_5_cse);
  assign nand_29_nl = ~(main_stage_v_1 & (~ mux_tmp_146));
  assign mux_168_nl = MUX_s_1_2_2((nand_29_nl), (mux_167_nl), or_1087_cse);
  assign IsZero_8U_23U_and_4_cse = core_wen & cfg_alu_algo_cfg_alu_algo_or_3_cse
      & (~ (mux_168_nl));
  assign IsZero_8U_23U_1_and_cse = chn_alu_out_and_8_cse & (~ or_dcpl_100);
  assign FpAdd_8U_23U_is_addition_and_cse = core_wen & (~ or_dcpl_100);
  assign nor_71_cse = ~(nor_269_cse | (cfg_precision!=2'b10) | cfg_alu_bypass_rsci_d
      | (~ chn_alu_in_rsci_bawt));
  assign and_489_cse = (~(or_937_cse & cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt)) & main_stage_v_1;
  assign and_231_rgt = and_dcpl_78 & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign and_233_rgt = and_dcpl_78 & or_dcpl_117 & (~ FpCmp_8U_23U_true_if_acc_4_itm_8);
  assign and_235_rgt = and_dcpl_78 & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign and_237_rgt = and_dcpl_78 & or_dcpl_119 & (~ FpCmp_8U_23U_true_if_acc_6_itm_8);
  assign and_239_rgt = and_dcpl_78 & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign and_241_rgt = and_dcpl_78 & or_dcpl_121 & (~ FpCmp_8U_23U_true_if_acc_8_itm_8);
  assign and_243_rgt = and_dcpl_78 & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign and_245_rgt = and_dcpl_78 & or_dcpl_123 & (~ FpCmp_8U_23U_true_if_acc_10_itm_8);
  assign nor_241_nl = ~((cfg_alu_algo_1_sva_st_23!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_4)
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5 | io_read_cfg_alu_bypass_rsc_svs_6
      | alu_loop_op_unequal_tmp_6);
  assign mux_176_nl = MUX_s_1_2_2(nor_264_cse, (nor_241_nl), FpAlu_8U_23U_equal_tmp_21);
  assign nor_243_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (FpAlu_8U_23U_equal_tmp_22
      & ((cfg_alu_algo_1_sva_st_24[0]) | (~((cfg_alu_algo_1_sva_st_24[1]) & FpAlu_8U_23U_nor_dfs_5)))));
  assign mux_177_nl = MUX_s_1_2_2((nor_243_nl), (mux_176_nl), or_1087_cse);
  assign IsNaN_8U_23U_aelse_and_12_cse = core_wen & (~ and_dcpl_32) & (mux_177_nl);
  assign FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse = (or_1087_cse & (~ alu_loop_op_unequal_tmp_6))
      | and_dcpl_165;
  assign mux_183_nl = MUX_s_1_2_2(or_tmp_305, or_tmp_395, or_1087_cse);
  assign or_426_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | or_tmp_305;
  assign mux_184_nl = MUX_s_1_2_2((or_426_nl), (mux_183_nl), or_tmp_402);
  assign AluOut_data_and_12_cse = core_wen & FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse
      & (~ (mux_184_nl));
  assign FpAlu_8U_23U_and_88_cse = core_wen & (~ and_dcpl_32) & (~ mux_tmp_171);
  assign or_441_nl = alu_loop_op_unequal_tmp_6 | or_tmp_416;
  assign mux_191_nl = MUX_s_1_2_2((or_441_nl), mux_tmp_171, FpAlu_8U_23U_equal_tmp_25);
  assign or_443_nl = (~ FpAlu_8U_23U_equal_tmp_25) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign mux_192_nl = MUX_s_1_2_2((or_443_nl), (mux_191_nl), FpAlu_8U_23U_equal_tmp_24);
  assign FpCmp_8U_23U_true_o_and_5_cse = core_wen & (~ and_dcpl_32) & (~ (mux_192_nl));
  assign mux_197_nl = MUX_s_1_2_2(or_tmp_269, or_tmp_395, or_1087_cse);
  assign or_453_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ FpAlu_8U_23U_equal_tmp_28) | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign nor_81_nl = ~(alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_equal_tmp_27));
  assign mux_198_nl = MUX_s_1_2_2((or_453_nl), (mux_197_nl), nor_81_nl);
  assign FpCmp_8U_23U_false_o_and_6_cse = core_wen & (~ and_dcpl_32) & (~ (mux_198_nl));
  assign nor_236_cse = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6);
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse = and_dcpl_165 | and_dcpl_168
      | and_dcpl_169;
  assign mux_201_nl = MUX_s_1_2_2(or_tmp_312, or_tmp_395, or_1087_cse);
  assign or_463_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ alu_loop_op_unequal_tmp_7) | io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign mux_202_nl = MUX_s_1_2_2((or_463_nl), (mux_201_nl), alu_loop_op_unequal_tmp_6);
  assign IntSaturation_33U_32U_and_11_cse = core_wen & (~ and_dcpl_32) & (~ (mux_202_nl));
  assign alu_loop_bypass_if_and_6_cse = (~ alu_loop_op_unequal_tmp_6) & and_dcpl_171;
  assign alu_loop_bypass_if_and_7_cse = alu_loop_op_unequal_tmp_6 & and_dcpl_171;
  assign AluOut_data_and_15_cse = core_wen & (and_dcpl_170 | alu_loop_bypass_if_and_6_cse
      | alu_loop_bypass_if_and_7_cse) & mux_tmp_53;
  assign and_485_nl = or_963_cse & (cfg_precision==2'b10) & main_stage_v_1 & cfg_alu_bypass_rsc_triosy_obj_bawt
      & cfg_alu_src_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt
      & (~ io_read_cfg_alu_bypass_rsc_svs_5);
  assign mux_213_nl = MUX_s_1_2_2((and_485_nl), and_484_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_214_nl = MUX_s_1_2_2(nor_197_cse, (mux_213_nl), or_1087_cse);
  assign FpAlu_8U_23U_and_94_cse = core_wen & (~ and_dcpl_32) & (mux_214_nl);
  assign mux_215_nl = MUX_s_1_2_2(or_381_cse, or_391_cse, and_489_cse);
  assign mux_216_nl = MUX_s_1_2_2(or_391_cse, (mux_215_nl), nor_71_cse);
  assign IsZero_8U_23U_and_6_cse = core_wen & (~ or_dcpl_109) & (~ (mux_216_nl));
  assign nor_208_nl = ~((cfg_precision!=2'b10) | (~ main_stage_v_1) | io_read_cfg_alu_bypass_rsc_svs_st_1
      | (~ cfg_alu_bypass_rsc_triosy_obj_bawt) | (~ cfg_alu_src_rsc_triosy_obj_bawt)
      | (~ cfg_alu_op_rsc_triosy_obj_bawt) | (~ cfg_alu_algo_rsc_triosy_obj_bawt)
      | io_read_cfg_alu_bypass_rsc_svs_5 | FpAlu_8U_23U_equal_tmp_1_mx0w0 | nor_202_cse);
  assign nor_210_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6 | (FpAlu_8U_23U_equal_tmp_21
      & ((cfg_alu_algo_1_sva_st_23[0]) | (~((cfg_alu_algo_1_sva_st_23[1]) & FpAlu_8U_23U_nor_dfs_4)))));
  assign mux_217_nl = MUX_s_1_2_2((nor_210_nl), (nor_208_nl), or_1087_cse);
  assign IsNaN_8U_23U_aelse_and_16_cse = core_wen & (~ and_dcpl_32) & (mux_217_nl);
  assign and_481_cse = or_963_cse & (cfg_precision==2'b10) & main_stage_v_1 & (~
      io_read_cfg_alu_bypass_rsc_svs_st_1) & cfg_alu_bypass_rsc_triosy_obj_bawt &
      cfg_alu_src_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt
      & (cfg_alu_algo_1_sva_2==2'b11) & (~ io_read_cfg_alu_bypass_rsc_svs_5);
  assign AluOut_data_and_5_cse = alu_loop_op_else_nor_dfs & and_dcpl_208;
  assign nor_204_nl = ~((cfg_precision[1]) | (~ or_963_cse));
  assign nor_390_nl = ~((~(FpAlu_8U_23U_equal_tmp_1_mx0w0 | (cfg_precision[0])))
      | io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_221_nl = MUX_s_1_2_2((nor_204_nl), or_963_cse, nor_390_nl);
  assign and_478_nl = main_stage_v_1 & cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt & (~ io_read_cfg_alu_bypass_rsc_svs_5)
      & (mux_221_nl);
  assign nor_205_nl = ~((~ or_tmp_402) | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6);
  assign mux_222_nl = MUX_s_1_2_2((nor_205_nl), (and_478_nl), or_1087_cse);
  assign AluOut_data_and_17_cse = core_wen & (~ and_dcpl_32) & (mux_222_nl);
  assign nor_202_cse = ~((~ cfg_alu_src_1_sva_st_1) | chn_alu_op_rsci_bawt);
  assign nor_201_cse = ~(nor_202_cse | (cfg_precision!=2'b10) | (~ main_stage_v_1)
      | io_read_cfg_alu_bypass_rsc_svs_st_1 | (~ cfg_alu_bypass_rsc_triosy_obj_bawt)
      | (~ cfg_alu_src_rsc_triosy_obj_bawt) | (~ cfg_alu_op_rsc_triosy_obj_bawt)
      | (~ cfg_alu_algo_rsc_triosy_obj_bawt) | (cfg_alu_algo_1_sva_2!=2'b00) | io_read_cfg_alu_bypass_rsc_svs_5);
  assign nor_200_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6
      | (~ FpAlu_8U_23U_equal_tmp_24));
  assign mux_224_nl = MUX_s_1_2_2((nor_200_nl), nor_201_cse, or_1087_cse);
  assign FpCmp_8U_23U_true_o_and_9_cse = core_wen & (~ and_dcpl_32) & (mux_224_nl);
  assign nor_197_cse = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6 |
      alu_loop_op_unequal_tmp_6);
  assign alu_loop_op_else_o_mux1h_1_itm = MUX_v_32_2_2(({1'b0 , (FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0[30:0])}),
      alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0, mux_337_itm);
  assign or_1050_cse = (cfg_precision!=2'b10);
  assign or_1055_cse = (cfg_alu_algo_1_sva_2!=2'b01);
  assign alu_loop_op_else_o_mux1h_3_itm = MUX_v_32_2_2(({1'b0 , (FpCmp_8U_23U_false_o_2_lpi_1_dfm_2[30:0])}),
      alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0, mux_337_itm);
  assign and_293_rgt = or_1087_cse & io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign alu_loop_op_else_o_mux1h_5_itm = MUX_v_32_2_2(({1'b0 , (FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0[30:0])}),
      alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0, mux_337_itm);
  assign alu_loop_op_else_o_mux1h_7_itm = MUX_v_32_2_2(({1'b0 , (FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0[30:0])}),
      alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0, mux_337_itm);
  assign IntSaturation_33U_32U_if_and_9_cse = core_wen & (~ and_dcpl_32) & not_tmp_232;
  assign mux_243_nl = MUX_s_1_2_2((~ mux_tmp_227), or_tmp_577, io_read_cfg_alu_bypass_rsc_svs_5);
  assign mux_244_nl = MUX_s_1_2_2(or_tmp_577, (~ mux_tmp_227), or_963_cse);
  assign mux_245_nl = MUX_s_1_2_2((mux_244_nl), or_tmp_577, io_read_cfg_alu_bypass_rsc_svs_5);
  assign mux_246_nl = MUX_s_1_2_2((mux_245_nl), (mux_243_nl), io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_247_nl = MUX_s_1_2_2(or_tmp_577, (mux_246_nl), main_stage_v_1);
  assign FpAlu_8U_23U_and_102_cse = core_wen & (~ and_dcpl_32) & (~ (mux_247_nl));
  assign FpAlu_8U_23U_or_cse = (alu_loop_op_else_nor_dfs & and_dcpl_214) | (FpAlu_8U_23U_equal_tmp_2_mx0w0
      & and_dcpl_214);
  assign and_297_m1c = (~ mux_tmp_323) & or_1087_cse;
  assign and_486_cse = cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse = and_dcpl_219 | and_dcpl_81 | and_dcpl_222
      | and_dcpl_225;
  assign mux_262_nl = MUX_s_1_2_2((~ mux_tmp_246), nand_tmp_20, and_451_cse);
  assign mux_263_nl = MUX_s_1_2_2((~ mux_tmp_246), nand_tmp_20, cfg_alu_algo_1_sva_st[0]);
  assign mux_264_nl = MUX_s_1_2_2((~ nand_tmp_20), mux_tmp_246, cfg_alu_algo_rsci_d[0]);
  assign mux_265_nl = MUX_s_1_2_2(mux_tmp_246, (~ nand_tmp_20), cfg_alu_algo_rsci_d[0]);
  assign mux_266_nl = MUX_s_1_2_2((mux_265_nl), (mux_264_nl), cfg_alu_algo_1_sva_st[0]);
  assign mux_267_nl = MUX_s_1_2_2((~ (mux_266_nl)), nand_tmp_20, cfg_alu_algo_rsci_d[1]);
  assign mux_268_nl = MUX_s_1_2_2((mux_267_nl), (mux_263_nl), cfg_alu_algo_1_sva_st[1]);
  assign mux_269_nl = MUX_s_1_2_2((mux_268_nl), (mux_262_nl), nor_6_cse);
  assign mux_270_nl = MUX_s_1_2_2(nand_tmp_20, (mux_269_nl), nor_5_cse);
  assign IsNaN_8U_23U_2_and_6_cse = core_wen & IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse
      & (~ (mux_270_nl));
  assign IsNaN_8U_23U_2_and_cse = core_wen & IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse;
  assign nor_177_cse = ~(and_486_cse | io_read_cfg_alu_bypass_rsc_svs_5);
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse = and_dcpl_222 | and_dcpl_227 | and_dcpl_229
      | and_dcpl_231;
  assign mux_281_cse = MUX_s_1_2_2(io_read_cfg_alu_bypass_rsc_svs_5, mux_tmp_265,
      and_486_cse);
  assign and_451_cse = (cfg_alu_algo_rsci_d==2'b11);
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse = and_dcpl_236 | and_dcpl_239 | and_dcpl_243;
  assign mux_306_nl = MUX_s_1_2_2(and_451_cse, and_tmp_35, and_489_cse);
  assign mux_307_nl = MUX_s_1_2_2(and_tmp_35, (mux_306_nl), nor_71_cse);
  assign IsNaN_8U_23U_2_and_9_cse = chn_alu_out_and_8_cse & IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse
      & (~ (mux_307_nl));
  assign mux_312_cse = MUX_s_1_2_2((~ (cfg_alu_algo_rsci_d[0])), (cfg_alu_algo_rsci_d[0]),
      cfg_alu_algo_rsci_d[1]);
  assign and_328_rgt = or_dcpl_14 & and_dcpl_234 & or_1087_cse & (~ (cfg_alu_algo_rsci_d[0]));
  assign FpAlu_8U_23U_mux1h_155_nl = MUX1HOT_s_1_5_2((reg_AluIn_data_sva_4_94_64_1_itm[0]),
      (FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1[0]), AluOut_data_2_0_sva_11, AluOut_data_2_0_lpi_1_dfm_3,
      (FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1[0]), {FpAlu_8U_23U_nor_dfs_6 , FpAlu_8U_23U_equal_tmp_26
      , FpAlu_8U_23U_equal_tmp_23 , FpAlu_8U_23U_and_30_cse , FpAlu_8U_23U_and_31_m1c});
  assign alu_loop_op_mux_204_mx1w1 = MUX_s_1_2_2((FpAlu_8U_23U_mux1h_155_nl), AluOut_data_1_0_sva_12,
      alu_loop_op_unequal_tmp_8);
  assign FpAlu_8U_23U_mux1h_154_nl = MUX1HOT_v_22_3_2((FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1[22:1]),
      AluOut_data_2_22_1_lpi_1_dfm_3, (FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1[22:1]),
      {FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_and_30_cse , FpAlu_8U_23U_and_31_m1c});
  assign FpAlu_8U_23U_not_22_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_and_11_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_mux1h_154_nl),
      (FpAlu_8U_23U_not_22_nl));
  assign AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0 = MUX1HOT_v_22_3_2((FpAlu_8U_23U_and_11_nl),
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4, (reg_AluIn_data_sva_4_94_64_1_itm[22:1]),
      {nor_437_cse , asn_267 , or_dcpl});
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13
      + 8'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl = nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl[7:0];
  assign FpAdd_8U_23U_and_31_nl = (~(FpAdd_8U_23U_and_2_tmp_3 | FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8))
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_19_nl = FpAdd_8U_23U_and_2_tmp_3 & (~ FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8)
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_32_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8 & FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_21_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_11)
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_mux1h_153_nl = MUX1HOT_v_8_7_2(FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13,
      (alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl), 8'b11111110, else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3,
      (FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1[30:23]), AluOut_data_2_30_23_lpi_1_dfm_3,
      (FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1[30:23]), {(FpAdd_8U_23U_and_31_nl)
      , (FpAdd_8U_23U_and_19_nl) , (FpAdd_8U_23U_and_32_nl) , (FpAdd_8U_23U_and_21_nl)
      , FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_and_30_cse , FpAlu_8U_23U_and_31_m1c});
  assign FpAlu_8U_23U_not_25_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_and_10_nl = MUX_v_8_2_2(8'b00000000, (FpAlu_8U_23U_mux1h_153_nl),
      (FpAlu_8U_23U_not_25_nl));
  assign nor_408_nl = ~(asn_267 | or_998_tmp);
  assign AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0 = MUX1HOT_v_8_3_2((FpAlu_8U_23U_and_10_nl),
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13, reg_AluIn_data_sva_4_94_64_itm, {(nor_408_nl)
      , asn_267 , or_998_tmp});
  assign or_16_cse = or_963_cse | io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign and_97_nl = (~((~(and_dcpl_4 & or_16_cse)) & main_stage_v_1)) & or_1050_cse
      & chn_alu_in_rsci_bawt & (~ cfg_alu_bypass_rsci_d) & or_1087_cse & (fsm_output[1]);
  assign alu_loop_op_2_Y_alu_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_97_nl);
  assign alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp = (AluIn_data_sva_127[30:23])
      == (else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23);
  assign alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp = (AluIn_data_sva_127[62:55])
      == (else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23);
  assign alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp = (AluIn_data_sva_127[94:87])
      == (else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23);
  assign alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp = (AluIn_data_sva_127[126:119])
      == (else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23);
  assign alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0
      = ~((AluIn_data_sva_127[127]) ^ (else_AluOp_data_3_lpi_1_dfm_mx0[31]));
  assign FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1)
      & alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp) | FpCmp_8U_23U_true_if_acc_10_itm_8;
  assign alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = (else_AluOp_data_3_lpi_1_dfm_mx0[30:0]!=31'b0000000000000000000000000000000);
  assign FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_4, FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_38_nl = ~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_4, (FpAdd_8U_23U_is_a_greater_oelse_not_38_nl));
  assign alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0
      = ~((AluIn_data_sva_127[95]) ^ (else_AluOp_data_2_lpi_1_dfm_mx0[31]));
  assign FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1)
      & alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp) | FpCmp_8U_23U_true_if_acc_8_itm_8;
  assign alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = (else_AluOp_data_2_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000)
      | (else_AluOp_data_2_lpi_1_dfm_mx3_30_0[30:23]!=8'b00000000);
  assign FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_5, FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_39_nl = ~ FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_5, (FpAdd_8U_23U_is_a_greater_oelse_not_39_nl));
  assign alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0
      = ~((AluIn_data_sva_127[63]) ^ (else_AluOp_data_1_lpi_1_dfm_mx0[31]));
  assign FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1)
      & alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp) | FpCmp_8U_23U_true_if_acc_6_itm_8;
  assign alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = (else_AluOp_data_1_lpi_1_dfm_mx2_30_0[22:0]!=23'b00000000000000000000000)
      | (else_AluOp_data_1_lpi_1_dfm_mx0[30:23]!=8'b00000000);
  assign FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_6, FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_40_nl = ~ FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_6, (FpAdd_8U_23U_is_a_greater_oelse_not_40_nl));
  assign alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0
      = ~((AluIn_data_sva_127[31]) ^ (else_AluOp_data_0_lpi_1_dfm_mx0[31]));
  assign FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1)
      & alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp) | FpCmp_8U_23U_true_if_acc_4_itm_8;
  assign alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = (else_AluOp_data_0_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000)
      | (else_AluOp_data_0_lpi_1_dfm_mx3_30_0[30:23]!=8'b00000000);
  assign FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_7, FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_41_nl = ~ FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0 = MUX_v_8_2_2(8'b00000000,
      z_out_7, (FpAdd_8U_23U_is_a_greater_oelse_not_41_nl));
  assign FpNormalize_8U_49U_if_or_itm_mx0w0 = (z_out_12[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign FpNormalize_8U_49U_if_or_1_itm_mx0w0 = (z_out_13[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign FpNormalize_8U_49U_if_or_2_itm_mx0w0 = (z_out_14[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign FpNormalize_8U_49U_if_or_3_itm_mx0w0 = (z_out_15[48:0]!=49'b0000000000000000000000000000000000000000000000000);
  assign FpAdd_8U_23U_and_4_tmp = (~ alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign FpNormalize_8U_49U_else_mux_4_nl = MUX_v_6_2_2((~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4),
      6'b1, FpAdd_8U_23U_if_3_if_and_tmp);
  assign nl_acc_nl = ({FpAdd_8U_23U_qr_2_lpi_1_dfm_7 , (~ FpAdd_8U_23U_if_3_if_and_tmp)})
      + conv_s2u_8_9({(~ FpAdd_8U_23U_if_3_if_and_tmp) , (FpNormalize_8U_49U_else_mux_4_nl)
      , 1'b1});
  assign acc_nl = nl_acc_nl[8:0];
  assign nor_436_nl = ~(FpAdd_8U_23U_and_4_tmp | mux_tmp);
  assign FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2(({{7{FpNormalize_8U_49U_oelse_not_9}},
      FpNormalize_8U_49U_oelse_not_9}), FpAdd_8U_23U_qr_2_lpi_1_dfm_7, (readslicef_9_8_1((acc_nl))),
      {(nor_436_nl) , FpAdd_8U_23U_and_4_tmp , mux_tmp});
  assign FpAdd_8U_23U_and_10_tmp = (~ alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1)
      & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign FpNormalize_8U_49U_else_mux_5_nl = MUX_v_6_2_2((~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5),
      6'b1, FpAdd_8U_23U_if_3_if_and_tmp_1);
  assign nl_acc_1_nl = ({FpAdd_8U_23U_qr_3_lpi_1_dfm_7 , (~ FpAdd_8U_23U_if_3_if_and_tmp_1)})
      + conv_s2u_8_9({(~ FpAdd_8U_23U_if_3_if_and_tmp_1) , (FpNormalize_8U_49U_else_mux_5_nl)
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[8:0];
  assign nor_435_nl = ~(FpAdd_8U_23U_and_10_tmp | mux_tmp_348);
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2(({{7{FpNormalize_8U_49U_oelse_not_11}},
      FpNormalize_8U_49U_oelse_not_11}), FpAdd_8U_23U_qr_3_lpi_1_dfm_7, (readslicef_9_8_1((acc_1_nl))),
      {(nor_435_nl) , FpAdd_8U_23U_and_10_tmp , mux_tmp_348});
  assign FpAdd_8U_23U_and_16_tmp = (~ alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1)
      & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign FpNormalize_8U_49U_else_mux_6_nl = MUX_v_6_2_2((~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6),
      6'b1, FpAdd_8U_23U_if_3_if_and_tmp_2);
  assign nl_acc_2_nl = ({FpAdd_8U_23U_qr_4_lpi_1_dfm_7 , (~ FpAdd_8U_23U_if_3_if_and_tmp_2)})
      + conv_s2u_8_9({(~ FpAdd_8U_23U_if_3_if_and_tmp_2) , (FpNormalize_8U_49U_else_mux_6_nl)
      , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[8:0];
  assign nor_434_nl = ~(FpAdd_8U_23U_and_16_tmp | mux_tmp_349);
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2(({{7{FpNormalize_8U_49U_oelse_not_13}},
      FpNormalize_8U_49U_oelse_not_13}), FpAdd_8U_23U_qr_4_lpi_1_dfm_7, (readslicef_9_8_1((acc_2_nl))),
      {(nor_434_nl) , FpAdd_8U_23U_and_16_tmp , mux_tmp_349});
  assign FpAdd_8U_23U_and_22_tmp = (~ alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1)
      & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign FpNormalize_8U_49U_else_mux_7_nl = MUX_v_6_2_2((~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7),
      6'b1, FpAdd_8U_23U_if_3_if_and_tmp_3);
  assign nl_acc_3_nl = ({FpAdd_8U_23U_qr_lpi_1_dfm_7 , (~ FpAdd_8U_23U_if_3_if_and_tmp_3)})
      + conv_s2u_8_9({(~ FpAdd_8U_23U_if_3_if_and_tmp_3) , (FpNormalize_8U_49U_else_mux_7_nl)
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[8:0];
  assign nor_433_nl = ~(FpAdd_8U_23U_and_22_tmp | mux_tmp_350);
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2(({{7{FpNormalize_8U_49U_oelse_not_15}},
      FpNormalize_8U_49U_oelse_not_15}), FpAdd_8U_23U_qr_lpi_1_dfm_7, (readslicef_9_8_1((acc_3_nl))),
      {(nor_433_nl) , FpAdd_8U_23U_and_22_tmp , mux_tmp_350});
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0 = nor_41_cse | (~ alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1);
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0 = nor_37_cse | (~ alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1);
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0 = nor_33_cse | (~ alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0 = nor_45_cse | (~ alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1);
  assign alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[126:96]!=31'b0000000000000000000000000000000);
  assign alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[94:64]!=31'b0000000000000000000000000000000);
  assign FpAlu_8U_23U_equal_tmp_1_mx0w0 = (cfg_alu_algo_1_sva_2==2'b11);
  assign alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = (chn_alu_in_rsci_d_mxwt[62:32]!=31'b0000000000000000000000000000000);
  assign IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_3_nor_10_tmp | (else_AluOp_data_3_lpi_1_dfm_mx0[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_3_nor_8_tmp | (else_AluOp_data_2_lpi_1_dfm_mx3_30_0[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_3_nor_6_tmp | (else_AluOp_data_1_lpi_1_dfm_mx0[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 = ~(IsNaN_8U_23U_3_nor_4_tmp | (else_AluOp_data_0_lpi_1_dfm_mx3_30_0[30:23]!=8'b11111111));
  assign FpAlu_8U_23U_o_0_sva_2_mx0w0 = (AluIn_data_sva_127[127:96]) != else_AluOp_data_3_lpi_1_dfm_mx0;
  assign AluOut_data_2_0_sva_3_mx0w0 = (AluIn_data_sva_127[95:64]) != else_AluOp_data_2_lpi_1_dfm_mx0;
  assign FpAlu_8U_23U_equal_tmp_mx0w0 = ~((cfg_alu_algo_1_sva_2!=2'b00));
  assign FpAlu_8U_23U_nor_dfs_mx0w0 = ~(FpAlu_8U_23U_equal_tmp_mx0w0 | FpAlu_8U_23U_equal_tmp_1_mx0w0
      | FpAlu_8U_23U_equal_tmp_2_mx0w0);
  assign FpAlu_8U_23U_equal_tmp_2_mx0w0 = (cfg_alu_algo_1_sva_2==2'b01);
  assign alu_loop_op_else_alu_loop_op_else_mux_3_nl = MUX_v_32_2_2((signext_32_31(alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0[31:1])),
      (alu_loop_op_else_else_else_else_ac_int_cctor_1_sva[32:1]), alu_loop_op_else_equal_tmp_2);
  assign alu_loop_op_else_not_18_nl = ~ FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (alu_loop_op_else_alu_loop_op_else_mux_3_nl), (alu_loop_op_else_not_18_nl));
  assign alu_loop_op_else_alu_loop_op_else_mux_2_nl = MUX_v_32_2_2((signext_32_31(alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0[31:1])),
      (alu_loop_op_else_else_else_else_ac_int_cctor_2_sva[32:1]), alu_loop_op_else_equal_tmp_2);
  assign alu_loop_op_else_not_20_nl = ~ FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (alu_loop_op_else_alu_loop_op_else_mux_2_nl), (alu_loop_op_else_not_20_nl));
  assign nl_alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl = conv_s2u_2_3(~ (alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0[31:30]))
      + 3'b1;
  assign alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl = nl_alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl[2:0];
  assign alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2 = readslicef_3_1_2((alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl));
  assign alu_loop_op_else_alu_loop_op_else_mux_1_nl = MUX_v_32_2_2((signext_32_31(alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0[31:1])),
      (alu_loop_op_else_else_else_else_ac_int_cctor_3_sva[32:1]), alu_loop_op_else_equal_tmp_2);
  assign alu_loop_op_else_not_22_nl = ~ FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (alu_loop_op_else_alu_loop_op_else_mux_1_nl), (alu_loop_op_else_not_22_nl));
  assign alu_loop_op_else_alu_loop_op_else_mux_nl = MUX_v_32_2_2((signext_32_31(alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0[31:1])),
      (alu_loop_op_else_else_else_else_ac_int_cctor_sva[32:1]), alu_loop_op_else_equal_tmp_2);
  assign alu_loop_op_else_not_21_nl = ~ FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (alu_loop_op_else_alu_loop_op_else_mux_nl), (alu_loop_op_else_not_21_nl));
  assign nl_alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl = conv_s2u_2_3(~ (alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0[31:30]))
      + 3'b1;
  assign alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl = nl_alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl[2:0];
  assign alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2 = readslicef_3_1_2((alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl));
  assign nl_alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl = conv_s2u_2_3(~ (alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0[31:30]))
      + 3'b1;
  assign alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl = nl_alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl[2:0];
  assign alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2 = readslicef_3_1_2((alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl));
  assign nl_alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl = conv_s2u_2_3(~ (alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0[31:30]))
      + 3'b1;
  assign alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl = nl_alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl[2:0];
  assign alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2 = readslicef_3_1_2((alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl));
  assign else_AluOp_data_3_lpi_1_dfm_mx0 = MUX_v_32_2_2(cfg_alu_op_1_sva_1, (chn_alu_op_rsci_d_mxwt[127:96]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23 = MUX_v_8_2_2((cfg_alu_op_1_sva_1[30:23]),
      (chn_alu_op_rsci_d_mxwt[126:119]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 = ~(IsNaN_8U_23U_2_nor_2_mx0w0
      | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2);
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 = ~((~((chn_alu_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[30:23]!=8'b11111111));
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 = ~((~((chn_alu_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000)))
      | (chn_alu_in_rsci_d_mxwt[62:55]!=8'b11111111));
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 = ~(IsNaN_8U_23U_2_nor_3_mx0w0
      | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2);
  assign alu_loop_op_else_nor_dfs = ~(FpAlu_8U_23U_equal_tmp_2_mx0w0 | FpAlu_8U_23U_equal_tmp_1_mx0w0
      | alu_loop_op_else_equal_tmp_2);
  assign alu_loop_op_else_equal_tmp_2 = (cfg_alu_algo_1_sva_2==2'b10);
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2 = ~((chn_alu_in_rsci_d_mxwt[126:119]==8'b11111111));
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2 = ~((chn_alu_in_rsci_d_mxwt[94:87]==8'b11111111));
  assign FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0 = (FpCmp_8U_23U_true_else_else_if_acc_4_itm_23
      & (~ FpCmp_8U_23U_false_else_if_acc_6_itm_8)) | FpCmp_8U_23U_true_if_acc_6_itm_8;
  assign FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0,
      FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2, or_dcpl_154);
  assign IsNaN_8U_23U_2_nor_3_mx0w0 = ~((chn_alu_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_2_nor_2_mx0w0 = ~((chn_alu_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000));
  assign alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2 = (chn_alu_in_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000);
  assign else_AluOp_data_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(cfg_alu_op_1_sva_1, (chn_alu_op_rsci_d_mxwt[31:0]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23 = MUX_v_8_2_2((cfg_alu_op_1_sva_1[30:23]),
      (chn_alu_op_rsci_d_mxwt[30:23]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_0_lpi_1_dfm_mx3_30_0 = MUX_v_31_2_2((cfg_alu_op_1_sva_1[30:0]),
      (chn_alu_op_rsci_d_mxwt[30:0]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_1_lpi_1_dfm_mx0 = MUX_v_32_2_2(cfg_alu_op_1_sva_1, (chn_alu_op_rsci_d_mxwt[63:32]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23 = MUX_v_8_2_2((cfg_alu_op_1_sva_1[30:23]),
      (chn_alu_op_rsci_d_mxwt[62:55]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_1_lpi_1_dfm_mx2_30_0 = MUX_v_31_2_2((cfg_alu_op_1_sva_1[30:0]),
      (chn_alu_op_rsci_d_mxwt[62:32]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_2_lpi_1_dfm_mx0 = MUX_v_32_2_2(cfg_alu_op_1_sva_1, (chn_alu_op_rsci_d_mxwt[95:64]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23 = MUX_v_8_2_2((cfg_alu_op_1_sva_1[30:23]),
      (chn_alu_op_rsci_d_mxwt[94:87]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_AluOp_data_2_lpi_1_dfm_mx3_30_0 = MUX_v_31_2_2((cfg_alu_op_1_sva_1[30:0]),
      (chn_alu_op_rsci_d_mxwt[94:64]), alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_19_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_1_sva, FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_1_sva,
      FpAdd_8U_23U_addend_larger_asn_19_mx0w1, FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_13_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_2_sva, FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_2_sva,
      FpAdd_8U_23U_addend_larger_asn_13_mx0w1, FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_7_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_3_sva, FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_3_sva,
      FpAdd_8U_23U_addend_larger_asn_7_mx0w1, FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_1_mx0w1,
      FpAdd_8U_23U_a_int_mant_p1_sva, FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6);
  assign FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_sva,
      FpAdd_8U_23U_addend_larger_asn_1_mx0w1, FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6);
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_qr_2_lpi_1_dfm_7[7:1])})
      + 8'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl = ({1'b1 , (FpAdd_8U_23U_qr_3_lpi_1_dfm_7[7:1])})
      + 8'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl = nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl[7:0];
  assign alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1 = readslicef_8_1_7((alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl));
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl = ({1'b1 , (FpAdd_8U_23U_qr_4_lpi_1_dfm_7[7:1])})
      + 8'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl = nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0];
  assign alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl));
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl = ({1'b1 , (FpAdd_8U_23U_qr_lpi_1_dfm_7[7:1])})
      + 8'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl = nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl[7:0];
  assign alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1 = readslicef_8_1_7((alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl));
  assign alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp = FpMantRNE_49U_24U_else_carry_sva
      & (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_sva = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_itm, FpNormalize_8U_49U_oelse_not_15);
  assign FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl),
      (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_3_sva
      & (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_3_sva = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_itm, FpNormalize_8U_49U_oelse_not_13);
  assign FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl),
      (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp = FpMantRNE_49U_24U_else_carry_2_sva
      & (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_2_sva = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_itm, FpNormalize_8U_49U_oelse_not_11);
  assign FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl),
      (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_1_sva
      & (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_1_sva = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm, FpNormalize_8U_49U_oelse_not_9);
  assign FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl),
      (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49:1]), FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign FpAlu_8U_23U_o_0_lpi_1_dfm_2 = MUX1HOT_s_1_5_2((reg_AluIn_data_sva_4_126_96_1_itm[0]),
      (FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1[0]), FpAlu_8U_23U_o_0_sva_9, FpAlu_8U_23U_o_0_lpi_1_dfm_4,
      (FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1[0]), {FpAlu_8U_23U_nor_dfs_6 , FpAlu_8U_23U_equal_tmp_26
      , FpAlu_8U_23U_equal_tmp_23 , FpAlu_8U_23U_and_44_cse , FpAlu_8U_23U_and_45_cse});
  assign FpAlu_8U_23U_mux1h_35_nl = MUX1HOT_v_22_4_2((reg_AluIn_data_sva_4_126_96_1_itm[22:1]),
      (FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1[22:1]), FpAlu_8U_23U_o_22_1_lpi_1_dfm_4,
      (FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1[22:1]), {FpAlu_8U_23U_nor_dfs_6 ,
      FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_and_44_cse , FpAlu_8U_23U_and_45_cse});
  assign FpAlu_8U_23U_not_21_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_o_22_1_lpi_1_dfm_2 = MUX_v_22_2_2(22'b0000000000000000000000,
      (FpAlu_8U_23U_mux1h_35_nl), (FpAlu_8U_23U_not_21_nl));
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl = FpAdd_8U_23U_o_expo_lpi_1_dfm_13
      + 8'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl = nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl[7:0];
  assign FpAdd_8U_23U_and_33_nl = (~(FpAdd_8U_23U_and_3_tmp_3 | FpAdd_8U_23U_is_inf_lpi_1_dfm_8))
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_25_nl = FpAdd_8U_23U_and_3_tmp_3 & (~ FpAdd_8U_23U_is_inf_lpi_1_dfm_8)
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_34_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm_8 & FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_27_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_lpi_1_dfm_11)
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_and_62_nl = IsNaN_8U_23U_land_lpi_1_dfm_11 & FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_mux1h_34_nl = MUX1HOT_v_8_8_2(FpAdd_8U_23U_o_expo_lpi_1_dfm_13,
      (alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl), 8'b11111110, else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3,
      reg_AluIn_data_sva_4_126_96_itm, (FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1[30:23]),
      FpAlu_8U_23U_o_30_23_lpi_1_dfm_4, (FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1[30:23]),
      {(FpAdd_8U_23U_and_33_nl) , (FpAdd_8U_23U_and_25_nl) , (FpAdd_8U_23U_and_34_nl)
      , (FpAdd_8U_23U_and_27_nl) , (FpAlu_8U_23U_and_62_nl) , FpAlu_8U_23U_equal_tmp_26
      , FpAlu_8U_23U_and_44_cse , FpAlu_8U_23U_and_45_cse});
  assign FpAlu_8U_23U_not_17_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_o_30_23_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000, (FpAlu_8U_23U_mux1h_34_nl),
      (FpAlu_8U_23U_not_17_nl));
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c = ~(IsNaN_8U_23U_1_land_lpi_1_dfm_9
      | IsNaN_8U_23U_land_lpi_1_dfm_11);
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c = ~(IsNaN_8U_23U_1_land_3_lpi_1_dfm_9
      | IsNaN_8U_23U_land_3_lpi_1_dfm_11);
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c = ~(IsNaN_8U_23U_1_land_2_lpi_1_dfm_9
      | IsNaN_8U_23U_land_2_lpi_1_dfm_11);
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c = ~(IsNaN_8U_23U_1_land_1_lpi_1_dfm_9
      | IsNaN_8U_23U_land_1_lpi_1_dfm_11);
  assign FpAlu_8U_23U_and_30_cse = (~ FpAlu_8U_23U_equal_tmp_32) & FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_31_m1c = FpAlu_8U_23U_equal_tmp_32 & FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_44_cse = (~ FpAlu_8U_23U_and_12_tmp) & FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_45_cse = FpAlu_8U_23U_and_12_tmp & FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_12_tmp = FpAlu_8U_23U_equal_tmp_35 & FpAlu_8U_23U_equal_tmp_32;
  assign main_stage_en_1 = chn_alu_in_rsci_bawt & (chn_alu_op_rsci_bawt | (~(cfg_alu_src_1_sva_st_1
      & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1))) & (cfg_alu_algo_rsc_triosy_obj_bawt
      | (~ main_stage_v_1)) & (cfg_alu_op_rsc_triosy_obj_bawt | (~ main_stage_v_1))
      & (cfg_alu_src_rsc_triosy_obj_bawt | (~ main_stage_v_1)) & (cfg_alu_bypass_rsc_triosy_obj_bawt
      | (~ main_stage_v_1)) & or_1087_cse;
  assign alu_loop_op_else_if_mux_8_nl = MUX_v_32_2_2(else_AluOp_data_0_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[31:0]), alu_loop_op_else_else_if_and_cse);
  assign alu_loop_op_else_if_mux_9_nl = MUX_v_32_2_2((~ (AluIn_data_sva_127[31:0])),
      (~ else_AluOp_data_0_lpi_1_dfm_mx0), alu_loop_op_else_else_if_and_cse);
  assign nl_acc_8_nl = conv_s2u_33_34({(alu_loop_op_else_if_mux_8_nl) , 1'b1}) +
      conv_s2u_33_34({(alu_loop_op_else_if_mux_9_nl) , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[33:0];
  assign alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0 = MUX_v_32_2_2(else_AluOp_data_0_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[31:0]), readslicef_34_1_33((acc_8_nl)));
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_1_sva = conv_s2s_32_33(AluIn_data_sva_127[31:0])
      + conv_s2s_32_33(else_AluOp_data_0_lpi_1_dfm_mx0);
  assign alu_loop_op_else_else_else_else_ac_int_cctor_1_sva = nl_alu_loop_op_else_else_else_else_ac_int_cctor_1_sva[32:0];
  assign alu_loop_op_else_if_mux_12_nl = MUX_v_32_2_2(else_AluOp_data_1_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[63:32]), alu_loop_op_else_else_if_and_cse);
  assign alu_loop_op_else_if_mux_13_nl = MUX_v_32_2_2((~ (AluIn_data_sva_127[63:32])),
      (~ else_AluOp_data_1_lpi_1_dfm_mx0), alu_loop_op_else_else_if_and_cse);
  assign nl_acc_10_nl = conv_s2u_33_34({(alu_loop_op_else_if_mux_12_nl) , 1'b1})
      + conv_s2u_33_34({(alu_loop_op_else_if_mux_13_nl) , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[33:0];
  assign alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0 = MUX_v_32_2_2(else_AluOp_data_1_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[63:32]), readslicef_34_1_33((acc_10_nl)));
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_2_sva = conv_s2s_32_33(AluIn_data_sva_127[63:32])
      + conv_s2s_32_33(else_AluOp_data_1_lpi_1_dfm_mx0);
  assign alu_loop_op_else_else_else_else_ac_int_cctor_2_sva = nl_alu_loop_op_else_else_else_else_ac_int_cctor_2_sva[32:0];
  assign alu_loop_op_else_if_mux_14_nl = MUX_v_32_2_2(else_AluOp_data_2_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[95:64]), alu_loop_op_else_else_if_and_1_cse);
  assign alu_loop_op_else_if_mux_15_nl = MUX_v_32_2_2((~ (AluIn_data_sva_127[95:64])),
      (~ else_AluOp_data_2_lpi_1_dfm_mx0), alu_loop_op_else_else_if_and_1_cse);
  assign nl_acc_11_nl = conv_s2u_33_34({(alu_loop_op_else_if_mux_14_nl) , 1'b1})
      + conv_s2u_33_34({(alu_loop_op_else_if_mux_15_nl) , 1'b1});
  assign acc_11_nl = nl_acc_11_nl[33:0];
  assign alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0 = MUX_v_32_2_2(else_AluOp_data_2_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[95:64]), readslicef_34_1_33((acc_11_nl)));
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_3_sva = conv_s2s_32_33(AluIn_data_sva_127[95:64])
      + conv_s2s_32_33(else_AluOp_data_2_lpi_1_dfm_mx0);
  assign alu_loop_op_else_else_else_else_ac_int_cctor_3_sva = nl_alu_loop_op_else_else_else_else_ac_int_cctor_3_sva[32:0];
  assign alu_loop_op_else_if_mux_10_nl = MUX_v_32_2_2(else_AluOp_data_3_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[127:96]), alu_loop_op_else_else_if_and_1_cse);
  assign alu_loop_op_else_if_mux_11_nl = MUX_v_32_2_2((~ (AluIn_data_sva_127[127:96])),
      (~ else_AluOp_data_3_lpi_1_dfm_mx0), alu_loop_op_else_else_if_and_1_cse);
  assign nl_acc_9_nl = conv_s2u_33_34({(alu_loop_op_else_if_mux_10_nl) , 1'b1}) +
      conv_s2u_33_34({(alu_loop_op_else_if_mux_11_nl) , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[33:0];
  assign alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(else_AluOp_data_3_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[127:96]), readslicef_34_1_33((acc_9_nl)));
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_sva = conv_s2s_32_33(AluIn_data_sva_127[127:96])
      + conv_s2s_32_33(else_AluOp_data_3_lpi_1_dfm_mx0);
  assign alu_loop_op_else_else_else_else_ac_int_cctor_sva = nl_alu_loop_op_else_else_else_else_ac_int_cctor_sva[32:0];
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl = nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7:0];
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1 = readslicef_8_1_7((alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl));
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl = nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0];
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = readslicef_8_1_7((alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl));
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl = nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7:0];
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1 = readslicef_8_1_7((alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl));
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl = ~(alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1
      | alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3);
  assign IntSaturation_33U_32U_and_3_nl = alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1
      & (~ alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3);
  assign IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1 = MUX1HOT_v_31_3_2(reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm,
      31'b1000000000000000000000000000000, 31'b111111111111111111111111111111, {(IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl)
      , (IntSaturation_33U_32U_and_3_nl) , alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3});
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl = ~(alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1
      | alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign IntSaturation_33U_32U_and_7_nl = alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1
      & (~ alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1 = MUX1HOT_v_31_3_2(reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm,
      31'b1000000000000000000000000000000, 31'b111111111111111111111111111111, {(IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl)
      , (IntSaturation_33U_32U_and_7_nl) , alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2});
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl = ~(alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1
      | alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2);
  assign IntSaturation_33U_32U_and_5_nl = alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1
      & (~ alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2);
  assign IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1 = MUX1HOT_v_31_3_2(reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm,
      31'b1000000000000000000000000000000, 31'b111111111111111111111111111111, {(IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl)
      , (IntSaturation_33U_32U_and_5_nl) , alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2});
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl = ~(alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1
      | alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2);
  assign IntSaturation_33U_32U_and_1_nl = alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1
      & (~ alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2);
  assign IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1 = MUX1HOT_v_31_3_2(reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm,
      31'b1000000000000000000000000000000, 31'b111111111111111111111111111111, {(IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl)
      , (IntSaturation_33U_32U_and_1_nl) , alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2});
  assign nl_alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl = conv_s2u_2_3({reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm
      , (reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm[30])}) + 3'b1;
  assign alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl = nl_alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl[2:0];
  assign alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1 = readslicef_3_1_2((alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl));
  assign nl_alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl = conv_s2u_2_3({reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm
      , (reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm[30])}) + 3'b1;
  assign alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl = nl_alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl[2:0];
  assign alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1 = readslicef_3_1_2((alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl));
  assign nl_alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl = conv_s2u_2_3({reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm
      , (reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm[30])}) + 3'b1;
  assign alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl = nl_alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl[2:0];
  assign alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1 = readslicef_3_1_2((alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl));
  assign nl_alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl = conv_s2u_2_3({reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm
      , (reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm[30])}) + 3'b1;
  assign alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl = nl_alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl[2:0];
  assign alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1 = readslicef_3_1_2((alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_4_nl = ({1'b1 , (AluIn_data_sva_127[30:23])})
      + conv_u2u_8_9(~ (else_AluOp_data_0_lpi_1_dfm_mx0[30:23])) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_4_nl = nl_FpCmp_8U_23U_false_else_if_acc_4_nl[8:0];
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_8_nl = ({1'b1 , (else_AluOp_data_0_lpi_1_dfm_mx3_30_0[22:0])})
      + conv_u2u_23_24(~ (AluIn_data_sva_127[22:0])) + 24'b1;
  assign FpCmp_8U_23U_true_else_else_if_acc_8_nl = nl_FpCmp_8U_23U_true_else_else_if_acc_8_nl[23:0];
  assign or_861_cse = (~((readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_4_nl)))
      | (~ (readslicef_24_1_23((FpCmp_8U_23U_true_else_else_if_acc_8_nl)))))) | FpCmp_8U_23U_true_if_acc_4_itm_8;
  assign nor_168_nl = ~((AluIn_data_sva_127[31]) | (~ or_tmp_668));
  assign and_446_nl = (else_mux_tmp_31_23[8]) & or_tmp_668;
  assign mux_339_nl = MUX_s_1_2_2((and_446_nl), (nor_168_nl), or_861_cse);
  assign asn_FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_nor_nl = ~((mux_339_nl) | IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2);
  assign FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0 = MUX_v_32_2_2((AluIn_data_sva_127[31:0]),
      else_AluOp_data_0_lpi_1_dfm_mx0, asn_FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_nor_nl);
  assign or_864_nl = (~(FpCmp_8U_23U_false_else_if_acc_6_itm_8 | (~ FpCmp_8U_23U_true_else_else_if_acc_4_itm_23)))
      | FpCmp_8U_23U_true_if_acc_6_itm_8;
  assign mux_340_nl = MUX_s_1_2_2((~ (else_mux_1_tmp_31_23[8])), (AluIn_data_sva_127[63]),
      or_864_nl);
  assign asn_FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_nor_nl = ~((~(((~ IsNaN_8U_23U_3_nor_6_tmp)
      & (else_mux_1_tmp_31_23[7:0]==8'b11111111)) | (mux_340_nl))) | IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1);
  assign FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0 = MUX_v_32_2_2((AluIn_data_sva_127[63:32]),
      else_AluOp_data_1_lpi_1_dfm_mx0, asn_FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_nor_nl);
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_7_nl = ({1'b1 , (else_AluOp_data_2_lpi_1_dfm_mx3_30_0[22:0])})
      + conv_u2u_23_24(~ (AluIn_data_sva_127[86:64])) + 24'b1;
  assign FpCmp_8U_23U_true_else_else_if_acc_7_nl = nl_FpCmp_8U_23U_true_else_else_if_acc_7_nl[23:0];
  assign nl_FpCmp_8U_23U_false_else_if_acc_8_nl = ({1'b1 , (AluIn_data_sva_127[94:87])})
      + conv_u2u_8_9(~ (else_AluOp_data_2_lpi_1_dfm_mx0[30:23])) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_8_nl = nl_FpCmp_8U_23U_false_else_if_acc_8_nl[8:0];
  assign or_867_cse = (~((~ (readslicef_24_1_23((FpCmp_8U_23U_true_else_else_if_acc_7_nl))))
      | (readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_8_nl))))) | FpCmp_8U_23U_true_if_acc_8_itm_8;
  assign nor_165_nl = ~((AluIn_data_sva_127[95]) | (~ or_tmp_674));
  assign and_444_nl = (else_mux_2_tmp_31_23[8]) & or_tmp_674;
  assign mux_341_nl = MUX_s_1_2_2((and_444_nl), (nor_165_nl), or_867_cse);
  assign asn_FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_nor_nl = ~((mux_341_nl) | IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1);
  assign FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0 = MUX_v_32_2_2((AluIn_data_sva_127[95:64]),
      else_AluOp_data_2_lpi_1_dfm_mx0, asn_FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_nor_nl);
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_6_nl = ({1'b1 , (else_AluOp_data_3_lpi_1_dfm_mx0[22:0])})
      + conv_u2u_23_24(~ (AluIn_data_sva_127[118:96])) + 24'b1;
  assign FpCmp_8U_23U_true_else_else_if_acc_6_nl = nl_FpCmp_8U_23U_true_else_else_if_acc_6_nl[23:0];
  assign nl_FpCmp_8U_23U_false_else_if_acc_10_nl = ({1'b1 , (AluIn_data_sva_127[126:119])})
      + conv_u2u_8_9(~ (else_AluOp_data_3_lpi_1_dfm_mx0[30:23])) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_10_nl = nl_FpCmp_8U_23U_false_else_if_acc_10_nl[8:0];
  assign or_871_cse = (~((~ (readslicef_24_1_23((FpCmp_8U_23U_true_else_else_if_acc_6_nl))))
      | (readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_10_nl))))) | FpCmp_8U_23U_true_if_acc_10_itm_8;
  assign nor_163_nl = ~((AluIn_data_sva_127[127]) | (~ or_tmp_678));
  assign and_443_nl = (else_mux_3_tmp_31_23[8]) & or_tmp_678;
  assign mux_342_nl = MUX_s_1_2_2((and_443_nl), (nor_163_nl), or_871_cse);
  assign asn_FpCmp_8U_23U_true_o_lpi_1_dfm_1_nor_nl = ~((mux_342_nl) | IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2);
  assign FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0 = MUX_v_32_2_2((AluIn_data_sva_127[127:96]),
      else_AluOp_data_3_lpi_1_dfm_mx0, asn_FpCmp_8U_23U_true_o_lpi_1_dfm_1_nor_nl);
  assign and_336_nl = (AluIn_data_sva_127[31]) & or_tmp_668;
  assign nor_162_nl = ~((else_mux_tmp_31_23[8]) | (~ or_tmp_668));
  assign mux_343_nl = MUX_s_1_2_2((nor_162_nl), (and_336_nl), or_861_cse);
  assign or_876_nl = (mux_343_nl) | IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
  assign FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0 = MUX_v_32_2_2(else_AluOp_data_0_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[31:0]), or_876_nl);
  assign and_338_nl = (AluIn_data_sva_127[95]) & or_tmp_674;
  assign nor_159_nl = ~((else_mux_2_tmp_31_23[8]) | (~ or_tmp_674));
  assign mux_344_nl = MUX_s_1_2_2((nor_159_nl), (and_338_nl), or_867_cse);
  assign or_880_nl = (mux_344_nl) | (~(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1
      | IsNaN_8U_23U_4_nor_2_itm_2));
  assign FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0 = MUX_v_32_2_2(else_AluOp_data_2_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[95:64]), or_880_nl);
  assign and_340_nl = (AluIn_data_sva_127[127]) & or_tmp_678;
  assign nor_156_nl = ~((else_mux_3_tmp_31_23[8]) | (~ or_tmp_678));
  assign mux_345_nl = MUX_s_1_2_2((nor_156_nl), (and_340_nl), or_871_cse);
  assign or_884_nl = (mux_345_nl) | (~(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1
      | IsNaN_8U_23U_4_nor_3_itm_3));
  assign FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0 = MUX_v_32_2_2(else_AluOp_data_3_lpi_1_dfm_mx0,
      (AluIn_data_sva_127[127:96]), or_884_nl);
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_nl = (~ FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0)
      & (else_AluOp_data_1_lpi_1_dfm_mx0[31]);
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_nl = FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0
      | (else_AluOp_data_1_lpi_1_dfm_mx0[31]);
  assign FpCmp_8U_23U_false_mux_4_nl = MUX_s_1_2_2((FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_nl),
      (FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_nl), AluIn_data_sva_127[63]);
  assign FpAlu_8U_23U_and_61_nl = ((FpCmp_8U_23U_false_mux_4_nl) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0)
      & (~ IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2) & FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpCmp_8U_23U_false_o_2_lpi_1_dfm_2 = MUX_v_32_2_2((AluIn_data_sva_127[63:32]),
      else_AluOp_data_1_lpi_1_dfm_mx0, FpAlu_8U_23U_and_61_nl);
  assign FpAlu_8U_23U_and_48_m1c = (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0) & FpAlu_8U_23U_and_34_m1c;
  assign FpAlu_8U_23U_and_34_m1c = (~ IsNaN_8U_23U_land_3_lpi_1_dfm_8) & FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_52_m1c = (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0) & FpAlu_8U_23U_and_36_m1c;
  assign FpAlu_8U_23U_and_36_m1c = (~ IsNaN_8U_23U_land_1_lpi_1_dfm_8) & FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_56_m1c = (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0) & FpAlu_8U_23U_and_38_m1c;
  assign FpAlu_8U_23U_and_38_m1c = (~ IsNaN_8U_23U_land_2_lpi_1_dfm_8) & FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_40_m1c = (~ IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0) & FpAlu_8U_23U_and_24_m1c;
  assign FpAlu_8U_23U_and_24_m1c = (~ IsNaN_8U_23U_land_lpi_1_dfm_8) & FpAlu_8U_23U_nor_dfs_mx0w0;
  assign nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_2_lpi_1_dfm_7)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4)
      + 9'b1;
  assign alu_loop_op_1_FpNormalize_8U_49U_acc_nl = nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_9 = FpNormalize_8U_49U_if_or_itm_2 & (readslicef_9_1_8((alu_loop_op_1_FpNormalize_8U_49U_acc_nl)));
  assign nl_alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_3_lpi_1_dfm_7)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5)
      + 9'b1;
  assign alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl = nl_alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_11 = FpNormalize_8U_49U_if_or_1_itm_2 & (readslicef_9_1_8((alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl)));
  assign nl_alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_4_lpi_1_dfm_7)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6)
      + 9'b1;
  assign alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl = nl_alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_13 = FpNormalize_8U_49U_if_or_2_itm_2 & (readslicef_9_1_8((alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl)));
  assign nl_alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl = ({1'b1 , (~ FpAdd_8U_23U_qr_lpi_1_dfm_7)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7)
      + 9'b1;
  assign alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl = nl_alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl[8:0];
  assign FpNormalize_8U_49U_oelse_not_15 = FpNormalize_8U_49U_if_or_3_itm_2 & (readslicef_9_1_8((alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl)));
  assign asn_267 = alu_loop_op_unequal_tmp_8 & (~ io_read_cfg_alu_bypass_rsc_svs_8);
  assign nl_FpCmp_8U_23U_true_if_acc_4_nl = ({1'b1 , else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23})
      + conv_u2u_8_9(~ (AluIn_data_sva_127[30:23])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_4_nl = nl_FpCmp_8U_23U_true_if_acc_4_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_4_itm_8 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_4_nl));
  assign IsNaN_8U_23U_3_nor_4_tmp = ~((else_AluOp_data_0_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000));
  assign nl_FpCmp_8U_23U_true_if_acc_6_nl = ({1'b1 , else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23})
      + conv_u2u_8_9(~ (AluIn_data_sva_127[62:55])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_6_nl = nl_FpCmp_8U_23U_true_if_acc_6_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_6_itm_8 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_6_nl));
  assign nl_FpCmp_8U_23U_false_else_if_acc_6_nl = ({1'b1 , (AluIn_data_sva_127[62:55])})
      + conv_u2u_8_9(~ (else_AluOp_data_1_lpi_1_dfm_mx2_30_0[30:23])) + 9'b1;
  assign FpCmp_8U_23U_false_else_if_acc_6_nl = nl_FpCmp_8U_23U_false_else_if_acc_6_nl[8:0];
  assign FpCmp_8U_23U_false_else_if_acc_6_itm_8 = readslicef_9_1_8((FpCmp_8U_23U_false_else_if_acc_6_nl));
  assign IsNaN_8U_23U_3_nor_6_tmp = ~((else_AluOp_data_1_lpi_1_dfm_mx2_30_0[22:0]!=23'b00000000000000000000000));
  assign else_else_mux_13_nl = MUX_v_23_2_2((cfg_alu_op_1_sva_1[22:0]), (chn_alu_op_rsci_d_mxwt[54:32]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_4_nl = ({1'b1 , (else_else_mux_13_nl)})
      + conv_u2u_23_24(~ (AluIn_data_sva_127[54:32])) + 24'b1;
  assign FpCmp_8U_23U_true_else_else_if_acc_4_nl = nl_FpCmp_8U_23U_true_else_else_if_acc_4_nl[23:0];
  assign FpCmp_8U_23U_true_else_else_if_acc_4_itm_23 = readslicef_24_1_23((FpCmp_8U_23U_true_else_else_if_acc_4_nl));
  assign nl_FpCmp_8U_23U_true_if_acc_8_nl = ({1'b1 , else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23})
      + conv_u2u_8_9(~ (AluIn_data_sva_127[94:87])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_8_nl = nl_FpCmp_8U_23U_true_if_acc_8_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_8_itm_8 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_8_nl));
  assign IsNaN_8U_23U_3_nor_8_tmp = ~((else_AluOp_data_2_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000));
  assign nl_FpCmp_8U_23U_true_if_acc_10_nl = ({1'b1 , else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23})
      + conv_u2u_8_9(~ (AluIn_data_sva_127[126:119])) + 9'b1;
  assign FpCmp_8U_23U_true_if_acc_10_nl = nl_FpCmp_8U_23U_true_if_acc_10_nl[8:0];
  assign FpCmp_8U_23U_true_if_acc_10_itm_8 = readslicef_9_1_8((FpCmp_8U_23U_true_if_acc_10_nl));
  assign IsNaN_8U_23U_3_nor_10_tmp = ~((else_AluOp_data_3_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000));
  assign else_mux_3_tmp_31_23 = MUX_v_9_2_2((cfg_alu_op_1_sva_1[31:23]), (chn_alu_op_rsci_d_mxwt[127:119]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_mux_2_tmp_31_23 = MUX_v_9_2_2((cfg_alu_op_1_sva_1[31:23]), (chn_alu_op_rsci_d_mxwt[95:87]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_mux_1_tmp_31_23 = MUX_v_9_2_2((cfg_alu_op_1_sva_1[31:23]), (chn_alu_op_rsci_d_mxwt[63:55]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign else_mux_tmp_31_23 = MUX_v_9_2_2((cfg_alu_op_1_sva_1[31:23]), (chn_alu_op_rsci_d_mxwt[31:23]),
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2);
  assign and_dcpl_2 = cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_dcpl_3 = cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt;
  assign and_dcpl_4 = and_dcpl_3 & and_dcpl_2;
  assign and_tmp = or_963_cse & cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt & or_1087_cse;
  assign or_tmp_9 = (~ main_stage_v_1) | io_read_cfg_alu_bypass_rsc_svs_st_1 | (cfg_alu_algo_1_sva_st_22!=2'b01)
      | (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01) | and_tmp;
  assign and_37_cse = cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt & or_1087_cse;
  assign or_967_nl = (~((cfg_alu_algo_1_sva_st_22!=2'b01) | (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01)))
      | and_tmp;
  assign mux_16_nl = MUX_s_1_2_2((or_967_nl), and_37_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_tmp_2 = MUX_s_1_2_2(or_1087_cse, (mux_16_nl), main_stage_v_1);
  assign or_tmp_15 = (~ main_stage_v_1) | io_read_cfg_alu_bypass_rsc_svs_st_1 | (cfg_alu_algo_1_sva_st_22!=2'b01)
      | and_tmp;
  assign or_965_nl = (~((cfg_alu_algo_1_sva_st_22!=2'b01))) | and_tmp;
  assign mux_24_nl = MUX_s_1_2_2((or_965_nl), and_37_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_tmp_10 = MUX_s_1_2_2(or_1087_cse, (mux_24_nl), main_stage_v_1);
  assign or_tmp_20 = (~ main_stage_v_1) | io_read_cfg_alu_bypass_rsc_svs_st_1 | and_tmp;
  assign nand_17_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_1 & (~(cfg_alu_bypass_rsc_triosy_obj_bawt
      & cfg_alu_src_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt
      & or_1087_cse)));
  assign mux_32_nl = MUX_s_1_2_2(or_1087_cse, (nand_17_nl), main_stage_v_1);
  assign mux_33_nl = MUX_s_1_2_2(or_tmp_20, (~ (mux_32_nl)), chn_alu_in_rsci_bawt);
  assign mux_34_itm = MUX_s_1_2_2((mux_33_nl), or_tmp_20, cfg_alu_bypass_rsci_d);
  assign not_tmp_24 = ~(cfg_alu_src_rsci_d & chn_alu_in_rsci_bawt);
  assign or_tmp_23 = nor_269_cse | cfg_alu_bypass_rsci_d | not_tmp_24;
  assign nor_371_nl = ~((~ main_stage_v_1) | io_read_cfg_alu_bypass_rsc_svs_st_1
      | (cfg_alu_algo_1_sva_st_22[0]) | (~((cfg_alu_algo_1_sva_st_22[1]) & cfg_alu_bypass_rsc_triosy_obj_bawt
      & cfg_alu_src_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt
      & or_963_cse)));
  assign nor_372_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign not_tmp_29 = MUX_s_1_2_2((nor_372_nl), (nor_371_nl), or_1087_cse);
  assign not_tmp_38 = ~((~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ main_stage_v_2));
  assign or_tmp_75 = (cfg_alu_algo_1_sva_st_24!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign nor_357_nl = ~((~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3));
  assign mux_56_nl = MUX_s_1_2_2((~ or_tmp_75), main_stage_v_2, or_1087_cse);
  assign or_87_nl = (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign not_tmp_57 = MUX_s_1_2_2((mux_56_nl), (nor_357_nl), or_87_nl);
  assign or_tmp_103 = io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_tmp_53 = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_1087_cse);
  assign or_tmp_218 = io_read_cfg_alu_bypass_rsc_svs_st_7 | alu_loop_op_unequal_tmp_8
      | io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign or_230_nl = nor_269_cse | FpAlu_8U_23U_equal_tmp_22 | alu_loop_op_unequal_tmp_7
      | io_read_cfg_alu_bypass_rsc_svs_7 | io_read_cfg_alu_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign or_233_nl = FpAlu_8U_23U_equal_tmp_22 | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_108_nl = MUX_s_1_2_2(or_tmp_218, (or_233_nl), or_1087_cse);
  assign mux_109_itm = MUX_s_1_2_2((mux_108_nl), (or_230_nl), FpAlu_8U_23U_equal_tmp_23);
  assign or_tmp_224 = io_read_cfg_alu_bypass_rsc_svs_st_7 | (~ main_stage_v_4);
  assign or_tmp_251 = alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign or_tmp_261 = (~ FpAlu_8U_23U_equal_tmp_31) | (~ FpAlu_8U_23U_equal_tmp_28)
      | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign or_tmp_269 = (~ FpAlu_8U_23U_equal_tmp_28) | alu_loop_op_unequal_tmp_7 |
      io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign or_tmp_280 = alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign or_tmp_293 = (~ FpAlu_8U_23U_equal_tmp_34) | (~ FpAlu_8U_23U_equal_tmp_31)
      | (~ FpAlu_8U_23U_equal_tmp_28) | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign or_tmp_305 = (~(FpAlu_8U_23U_equal_tmp_22 | alu_loop_op_unequal_tmp_7))
      | io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign or_tmp_309 = (~ alu_loop_op_unequal_tmp_8) | io_read_cfg_alu_bypass_rsc_svs_8
      | (~ main_stage_v_4);
  assign or_323_nl = io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_141_nl = MUX_s_1_2_2((or_323_nl), or_tmp_305, or_1087_cse);
  assign mux_142_nl = MUX_s_1_2_2(or_tmp_309, or_tmp_305, or_1087_cse);
  assign mux_143_itm = MUX_s_1_2_2((mux_142_nl), (mux_141_nl), FpAlu_8U_23U_equal_tmp_23);
  assign or_tmp_312 = (~ alu_loop_op_unequal_tmp_7) | io_read_cfg_alu_bypass_rsc_svs_7
      | (~ main_stage_v_3);
  assign or_tmp_315 = nor_269_cse | (cfg_alu_algo_1_sva_st_24!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3) | (cfg_precision!=2'b10);
  assign or_tmp_347 = nor_269_cse | (~ main_stage_v_2) | (cfg_precision!=2'b10);
  assign not_tmp_152 = ~((cfg_alu_algo_1_sva_st_22!=2'b10));
  assign or_386_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 | (cfg_alu_algo_1_sva_st_22!=2'b10);
  assign nor_248_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_1 | not_tmp_152);
  assign mux_tmp_146 = MUX_s_1_2_2((nor_248_nl), (or_386_nl), io_read_cfg_alu_bypass_rsc_svs_5);
  assign or_383_nl = (~ cfg_alu_src_1_sva_st_1) | chn_alu_op_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_1
      | (cfg_alu_algo_1_sva_st_22!=2'b10);
  assign mux_162_nl = MUX_s_1_2_2(mux_tmp_146, (or_383_nl), and_486_cse);
  assign nand_tmp_13 = ~(main_stage_v_1 & (~ (mux_162_nl)));
  assign nor_379_nl = ~((~ cfg_alu_src_1_sva_st_1) | chn_alu_op_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_1
      | not_tmp_152);
  assign mux_163_nl = MUX_s_1_2_2(mux_tmp_146, (nor_379_nl), and_486_cse);
  assign not_tmp_157 = main_stage_v_1 & (mux_163_nl);
  assign or_391_cse = (cfg_alu_algo_1_sva_st!=2'b10);
  assign or_381_cse = (cfg_alu_algo_rsci_d!=2'b10);
  assign or_tmp_382 = (cfg_alu_algo_1_sva_st!=2'b01);
  assign or_tmp_386 = cfg_alu_bypass_rsci_d | (~ chn_alu_in_rsci_bawt);
  assign nor_tmp_74 = io_read_cfg_alu_bypass_rsc_svs_5 & io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign or_tmp_395 = io_read_cfg_alu_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign or_417_nl = io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign or_419_nl = io_read_cfg_alu_bypass_rsc_svs_7 | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_178_nl = MUX_s_1_2_2((or_419_nl), (or_417_nl), alu_loop_op_unequal_tmp_7);
  assign mux_tmp_164 = MUX_s_1_2_2(or_tmp_312, (mux_178_nl), FpAlu_8U_23U_equal_tmp_22);
  assign mux_tmp_165 = MUX_s_1_2_2(mux_tmp_164, or_tmp_395, or_1087_cse);
  assign or_tmp_402 = alu_loop_op_unequal_tmp_6 | FpAlu_8U_23U_equal_tmp_21;
  assign or_428_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign mux_185_nl = MUX_s_1_2_2(or_tmp_251, or_tmp_395, or_1087_cse);
  assign mux_tmp_171 = MUX_s_1_2_2((mux_185_nl), (or_428_nl), alu_loop_op_unequal_tmp_6);
  assign or_tmp_409 = alu_loop_op_unequal_tmp_6 | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_432_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7 | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_187_nl = MUX_s_1_2_2(or_tmp_280, or_tmp_395, or_1087_cse);
  assign mux_tmp_173 = MUX_s_1_2_2((mux_187_nl), (or_432_nl), or_tmp_409);
  assign or_tmp_416 = nor_269_cse | io_read_cfg_alu_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign and_484_cse = main_stage_v_1 & cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt & (~ io_read_cfg_alu_bypass_rsc_svs_5);
  assign and_474_nl = or_963_cse & or_1050_cse & main_stage_v_1 & cfg_alu_bypass_rsc_triosy_obj_bawt
      & cfg_alu_src_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt
      & (~ io_read_cfg_alu_bypass_rsc_svs_5);
  assign mux_233_nl = MUX_s_1_2_2((and_474_nl), and_484_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nor_187_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6 | (~
      alu_loop_op_unequal_tmp_6));
  assign not_tmp_232 = MUX_s_1_2_2((nor_187_nl), (mux_233_nl), or_1087_cse);
  assign or_tmp_577 = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | io_read_cfg_alu_bypass_rsc_svs_6 | (~ main_stage_v_2);
  assign mux_tmp_227 = MUX_s_1_2_2((~ or_tmp_395), and_dcpl_4, or_1087_cse);
  assign or_tmp_583 = (cfg_alu_algo_1_sva_st_22[0]) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt;
  assign or_tmp_585 = (~ (cfg_alu_algo_1_sva_st_22[0])) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt;
  assign mux_251_nl = MUX_s_1_2_2((cfg_alu_algo_1_sva_st_22[0]), (~ (cfg_alu_algo_1_sva_st_22[0])),
      cfg_alu_algo_1_sva_2[0]);
  assign or_609_nl = io_read_cfg_alu_bypass_rsc_svs_5 | (cfg_alu_algo_1_sva_2[1])
      | (mux_251_nl);
  assign mux_tmp_237 = MUX_s_1_2_2((or_609_nl), (cfg_alu_algo_1_sva_st_22[0]), cfg_alu_algo_1_sva_st_22[1]);
  assign or_601_nl = io_read_cfg_alu_bypass_rsc_svs_5 | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt;
  assign mux_248_nl = MUX_s_1_2_2(io_read_cfg_alu_bypass_rsc_svs_5, (or_601_nl),
      and_486_cse);
  assign mux_249_nl = MUX_s_1_2_2(or_tmp_583, or_tmp_585, cfg_alu_algo_1_sva_2[0]);
  assign or_607_nl = io_read_cfg_alu_bypass_rsc_svs_5 | (cfg_alu_algo_1_sva_2[1])
      | (mux_249_nl);
  assign mux_250_nl = MUX_s_1_2_2((or_607_nl), or_tmp_583, cfg_alu_algo_1_sva_st_22[1]);
  assign mux_253_nl = MUX_s_1_2_2(mux_tmp_237, (mux_250_nl), and_501_cse);
  assign mux_254_nl = MUX_s_1_2_2((mux_253_nl), (mux_248_nl), io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nand_tmp_20 = ~(main_stage_v_1 & (~ (mux_254_nl)));
  assign or_610_nl = (~ io_read_cfg_alu_bypass_rsc_svs_5) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt;
  assign mux_255_nl = MUX_s_1_2_2((~ io_read_cfg_alu_bypass_rsc_svs_5), (or_610_nl),
      and_486_cse);
  assign mux_256_nl = MUX_s_1_2_2(or_tmp_585, or_tmp_583, cfg_alu_algo_1_sva_2[0]);
  assign or_612_nl = io_read_cfg_alu_bypass_rsc_svs_5 | (cfg_alu_algo_1_sva_2[1]);
  assign mux_257_nl = MUX_s_1_2_2((mux_256_nl), or_1087_cse, or_612_nl);
  assign mux_258_nl = MUX_s_1_2_2((mux_257_nl), or_tmp_585, cfg_alu_algo_1_sva_st_22[1]);
  assign mux_259_nl = MUX_s_1_2_2((~ mux_tmp_237), (mux_258_nl), and_501_cse);
  assign mux_260_nl = MUX_s_1_2_2((mux_259_nl), (mux_255_nl), io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_tmp_246 = MUX_s_1_2_2(or_1087_cse, (mux_260_nl), main_stage_v_1);
  assign not_tmp_259 = ~((cfg_alu_algo_1_sva_st[0]) & ((cfg_alu_algo_1_sva_st_20!=2'b01)));
  assign or_tmp_596 = nor_71_cse | (cfg_alu_algo_1_sva_st[1]) | not_tmp_259;
  assign or_tmp_597 = (cfg_alu_algo_1_sva_st[1]) | not_tmp_259;
  assign not_tmp_261 = ~((reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01) | (~ or_tmp_597));
  assign or_629_nl = (~ (cfg_alu_algo_1_sva_st[0])) | (cfg_alu_algo_1_sva_st_20!=2'b01)
      | (cfg_alu_algo_rsci_d!=2'b01);
  assign mux_279_nl = MUX_s_1_2_2((or_629_nl), (cfg_alu_algo_1_sva_st[0]), cfg_alu_algo_1_sva_st[1]);
  assign mux_tmp_265 = MUX_s_1_2_2((mux_279_nl), mux_312_cse, nor_6_cse);
  assign mux_282_cse = MUX_s_1_2_2((~ (cfg_alu_algo_1_sva_st_22[1])), (cfg_alu_algo_1_sva_st_22[1]),
      cfg_alu_algo_1_sva_st_22[0]);
  assign or_632_cse = (cfg_alu_algo_1_sva_st_22!=2'b10);
  assign nor_117_nl = ~(io_read_cfg_alu_bypass_rsc_svs_5 | (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01)
      | (cfg_alu_algo_1_sva_st_28!=2'b01) | (cfg_alu_algo_1_sva_2!=2'b01));
  assign mux_tmp_268 = MUX_s_1_2_2(or_632_cse, mux_282_cse, nor_117_nl);
  assign nor_124_nl = ~(io_read_cfg_alu_bypass_rsc_svs_5 | (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01)
      | (cfg_alu_algo_1_sva_2!=2'b01));
  assign mux_tmp_281 = MUX_s_1_2_2(or_632_cse, mux_282_cse, nor_124_nl);
  assign nor_tmp_126 = (cfg_alu_algo_1_sva_st==2'b11);
  assign and_tmp_35 = (cfg_alu_algo_1_sva_st[0]) & or_28_cse;
  assign mux_310_nl = MUX_s_1_2_2((~ (cfg_alu_algo_1_sva_st[0])), (cfg_alu_algo_1_sva_st[0]),
      cfg_alu_algo_1_sva_st[1]);
  assign nor_143_nl = ~((cfg_alu_algo_1_sva_st_20!=2'b01));
  assign mux_tmp_296 = MUX_s_1_2_2(or_391_cse, (mux_310_nl), nor_143_nl);
  assign or_dcpl_14 = ~((~(and_dcpl_3 & and_dcpl_2 & or_16_cse)) & main_stage_v_1);
  assign and_dcpl_28 = and_dcpl_3 & cfg_alu_op_rsc_triosy_obj_bawt;
  assign and_dcpl_30 = (~((~(and_dcpl_28 & (chn_alu_op_rsci_bawt | io_read_cfg_alu_bypass_rsc_svs_st_1)
      & cfg_alu_algo_rsc_triosy_obj_bawt)) & main_stage_v_1)) & or_1087_cse;
  assign and_dcpl_32 = (~ chn_alu_out_rsci_bawt) & reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_33 = (~ chn_alu_op_rsci_bawt) & cfg_alu_src_1_sva_st_1;
  assign and_dcpl_34 = and_dcpl_33 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign or_dcpl_20 = ~(cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt);
  assign and_dcpl_35 = (or_dcpl_20 | and_dcpl_34) & main_stage_v_1;
  assign and_dcpl_37 = main_stage_v_4 & io_read_cfg_alu_bypass_rsc_svs_8;
  assign and_dcpl_40 = main_stage_v_4 & (~ io_read_cfg_alu_bypass_rsc_svs_8) & or_1087_cse;
  assign or_dcpl_23 = and_dcpl_32 | (~ main_stage_v_4);
  assign and_dcpl_43 = or_1087_cse & main_stage_v_4;
  assign and_dcpl_45 = (~ main_stage_v_4) & chn_alu_out_rsci_bawt & reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_46 = chn_alu_in_rsci_bawt & (~ cfg_alu_bypass_rsci_d);
  assign and_dcpl_53 = cfg_alu_src_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt
      & cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_dcpl_64 = or_16_cse & or_1087_cse & and_dcpl_28 & cfg_alu_algo_rsc_triosy_obj_bawt
      & main_stage_v_1;
  assign and_dcpl_70 = and_dcpl_28 & or_1087_cse;
  assign or_dcpl_46 = or_1050_cse | and_dcpl_32;
  assign or_dcpl_49 = and_dcpl_35 | and_dcpl_32;
  assign and_dcpl_77 = (cfg_precision==2'b10);
  assign and_dcpl_78 = and_dcpl_77 & or_1087_cse;
  assign and_dcpl_80 = or_dcpl_14 & or_1050_cse;
  assign and_dcpl_81 = and_dcpl_80 & or_1087_cse;
  assign and_dcpl_83 = or_dcpl_14 & and_dcpl_46 & or_1087_cse;
  assign and_dcpl_89 = chn_alu_in_rsci_bawt & cfg_alu_bypass_rsci_d;
  assign and_dcpl_96 = or_1087_cse & main_stage_v_2;
  assign and_dcpl_99 = or_1050_cse & or_1087_cse;
  assign and_dcpl_108 = or_1087_cse & alu_loop_op_unequal_tmp_7;
  assign or_tmp_657 = (~ or_1087_cse) | io_read_cfg_alu_bypass_rsc_svs_7;
  assign mux_tmp_311 = MUX_s_1_2_2(io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_7,
      or_1087_cse);
  assign nor_tmp_144 = alu_loop_op_unequal_tmp_7 & main_stage_v_3;
  assign and_dcpl_127 = nor_tmp_144 & or_1087_cse;
  assign or_dcpl_85 = or_1050_cse | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | and_dcpl_32;
  assign or_dcpl_86 = (cfg_alu_algo_1_sva_st_23!=2'b10);
  assign or_dcpl_89 = or_dcpl_46 | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_dcpl_86;
  assign or_dcpl_91 = or_1050_cse | (~ main_stage_v_2);
  assign or_dcpl_100 = or_dcpl_20 | and_dcpl_32 | (cfg_precision!=2'b10) | (cfg_alu_algo_1_sva_st_22[0])
      | and_dcpl_33 | (~ (cfg_alu_algo_1_sva_st_22[1])) | io_read_cfg_alu_bypass_rsc_svs_st_1
      | (~ main_stage_v_1);
  assign or_dcpl_109 = and_dcpl_35 | or_tmp_386 | (~ (cfg_precision[1])) | and_dcpl_32
      | (cfg_precision[0]);
  assign or_dcpl_117 = (~ alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1;
  assign or_dcpl_119 = (~ alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1;
  assign or_dcpl_121 = (~ alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1;
  assign or_dcpl_123 = (~ alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp)
      | FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1;
  assign and_dcpl_165 = or_1087_cse & alu_loop_op_unequal_tmp_6;
  assign and_dcpl_167 = or_1087_cse & (cfg_precision[1]);
  assign and_dcpl_168 = and_dcpl_167 & (~ (cfg_precision[0])) & (~ alu_loop_op_unequal_tmp_6);
  assign and_dcpl_169 = and_dcpl_99 & (~ alu_loop_op_unequal_tmp_6);
  assign and_dcpl_170 = or_1087_cse & io_read_cfg_alu_bypass_rsc_svs_6;
  assign and_dcpl_171 = or_1087_cse & (~ io_read_cfg_alu_bypass_rsc_svs_6);
  assign or_dcpl_125 = io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ (cfg_alu_algo_1_sva_st_23[1]));
  assign or_dcpl_127 = or_dcpl_91 | and_dcpl_32;
  assign and_dcpl_175 = ~((cfg_precision[0]) | (cfg_alu_algo_1_sva_st_22!=2'b10)
      | io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign and_dcpl_179 = and_dcpl_70 & cfg_alu_algo_rsc_triosy_obj_bawt & (cfg_precision[1])
      & or_963_cse;
  assign and_dcpl_207 = and_dcpl_167 & (~ (cfg_precision[0])) & (~ io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign and_dcpl_208 = (or_1050_cse | io_read_cfg_alu_bypass_rsc_svs_st_1) & or_1087_cse;
  assign mux_337_itm = MUX_s_1_2_2(and_dcpl_99, or_dcpl_46, alu_loop_op_unequal_tmp_6);
  assign mux_tmp_323 = ~(io_read_cfg_alu_bypass_rsc_svs_st_1 | and_dcpl_77);
  assign and_dcpl_214 = mux_tmp_323 & or_1087_cse;
  assign and_dcpl_217 = and_dcpl_77 & (~ (cfg_alu_algo_rsci_d[0]));
  assign and_dcpl_219 = or_dcpl_14 & and_dcpl_217 & or_1087_cse & (~ (cfg_alu_algo_rsci_d[1]));
  assign and_dcpl_222 = or_dcpl_14 & and_dcpl_77 & (cfg_alu_algo_rsci_d[0]) & or_1087_cse;
  assign and_dcpl_225 = or_dcpl_14 & and_dcpl_217 & or_1087_cse & (cfg_alu_algo_rsci_d[1]);
  assign or_dcpl_154 = (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01);
  assign and_dcpl_227 = and_dcpl_80 & or_1087_cse & (~ (cfg_alu_algo_1_sva_st[1]));
  assign and_dcpl_229 = or_dcpl_14 & and_dcpl_217 & or_1087_cse;
  assign and_dcpl_231 = and_dcpl_80 & or_1087_cse & (cfg_alu_algo_1_sva_st[1]);
  assign and_dcpl_234 = and_dcpl_46 & and_dcpl_77;
  assign and_dcpl_236 = or_dcpl_14 & and_dcpl_234 & (cfg_alu_algo_rsci_d==2'b00)
      & or_1087_cse;
  assign and_dcpl_239 = or_dcpl_14 & and_dcpl_234 & or_1087_cse & (cfg_alu_algo_rsci_d[0]);
  assign and_dcpl_243 = or_dcpl_14 & and_dcpl_234 & (cfg_alu_algo_rsci_d==2'b10)
      & or_1087_cse;
  assign or_tmp_668 = IsNaN_8U_23U_3_nor_4_tmp | (else_mux_tmp_31_23[7:0]!=8'b11111111);
  assign or_tmp_674 = IsNaN_8U_23U_3_nor_8_tmp | (else_mux_2_tmp_31_23[7:0]!=8'b11111111);
  assign or_tmp_678 = IsNaN_8U_23U_3_nor_10_tmp | (else_mux_3_tmp_31_23[7:0]!=8'b11111111);
  assign or_tmp_695 = or_dcpl_14 & or_1087_cse & chn_alu_in_rsci_bawt & (fsm_output[1]);
  assign and_357_cse = or_dcpl_14 & or_1087_cse & and_dcpl_46 & cfg_alu_src_rsci_d
      & (fsm_output[1]);
  assign chn_alu_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign chn_alu_op_rsci_ld_core_psct_mx0c1 = or_1087_cse & cfg_alu_bypass_rsc_triosy_obj_bawt
      & chn_alu_op_rsci_bawt & cfg_alu_src_1_sva_st_1 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1)
      & main_stage_v_1 & and_dcpl_53 & (or_tmp_386 | (~ cfg_alu_src_rsci_d));
  assign main_stage_v_1_mx0c1 = or_1087_cse & cfg_alu_bypass_rsc_triosy_obj_bawt
      & or_16_cse & and_dcpl_53 & (~ chn_alu_in_rsci_bawt) & main_stage_v_1;
  assign cfg_alu_src_1_sva_st_1_mx0c1 = (or_dcpl_14 & and_dcpl_89 & or_1087_cse &
      (fsm_output[1])) | (and_dcpl_30 & and_dcpl_89 & cfg_alu_src_1_sva_st_1);
  assign main_stage_v_2_mx0c1 = (or_dcpl_20 | and_dcpl_34 | (~ main_stage_v_1)) &
      and_dcpl_96;
  assign main_stage_v_3_mx0c1 = main_stage_v_3 & (~ main_stage_v_2) & or_1087_cse;
  assign main_stage_v_4_mx0c1 = (~ main_stage_v_3) & main_stage_v_4 & or_1087_cse;
  assign FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1 = and_dcpl_179 & and_dcpl_175 & main_stage_v_1
      & (~ FpCmp_8U_23U_true_if_acc_4_itm_8) & or_dcpl_117;
  assign FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1 = and_dcpl_179 & and_dcpl_175 & main_stage_v_1
      & (~ FpCmp_8U_23U_true_if_acc_6_itm_8) & or_dcpl_119;
  assign FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1 = and_dcpl_179 & and_dcpl_175 & main_stage_v_1
      & (~ FpCmp_8U_23U_true_if_acc_8_itm_8) & or_dcpl_121;
  assign FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1 = and_dcpl_179 & and_dcpl_175 & main_stage_v_1
      & (~ FpCmp_8U_23U_true_if_acc_10_itm_8) & or_dcpl_123;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = ({1'b1 , (AluIn_data_sva_127[22:0])})
      + conv_u2u_23_24(~ (else_AluOp_data_0_lpi_1_dfm_mx0[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , (AluIn_data_sva_127[54:32])})
      + conv_u2u_23_24(~ (else_AluOp_data_1_lpi_1_dfm_mx0[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , (AluIn_data_sva_127[86:64])})
      + conv_u2u_23_24(~ (else_AluOp_data_2_lpi_1_dfm_mx0[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , (AluIn_data_sva_127[118:96])})
      + conv_u2u_23_24(~ (else_AluOp_data_3_lpi_1_dfm_mx0[22:0])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23:0];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl));
  assign chn_alu_in_rsci_oswt_unreg = or_tmp_695;
  assign chn_alu_op_rsci_oswt_unreg = and_dcpl_70 & cfg_alu_algo_rsc_triosy_obj_bawt
      & chn_alu_op_rsci_bawt & cfg_alu_src_1_sva_st_1 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1)
      & main_stage_v_1;
  assign chn_alu_out_rsci_oswt_unreg = chn_alu_out_rsci_bawt & reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff = and_dcpl_64;
  assign and_dcpl_269 = nor_397_cse & (~ FpAlu_8U_23U_equal_tmp_23);
  assign or_996_tmp = (and_dcpl_269 & FpAlu_8U_23U_nor_dfs_6 & IsNaN_8U_23U_land_1_lpi_1_dfm_11)
      | io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_997_tmp = (and_dcpl_269 & FpAlu_8U_23U_nor_dfs_6 & IsNaN_8U_23U_land_2_lpi_1_dfm_11)
      | io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_998_tmp = (and_dcpl_269 & IsNaN_8U_23U_land_3_lpi_1_dfm_11 & FpAlu_8U_23U_nor_dfs_6)
      | io_read_cfg_alu_bypass_rsc_svs_8;
  assign and_dcpl = core_wen & main_stage_v_3;
  assign and_dcpl_349 = cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt;
  assign FpAdd_8U_23U_if_3_if_and_tmp = (fsm_output[1]) & (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_if_3_if_and_tmp_1 = (fsm_output[1]) & (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_if_3_if_and_tmp_2 = (fsm_output[1]) & (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_if_3_if_and_tmp_3 = (fsm_output[1]) & (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp = (fsm_output[1]) & (~((~(FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1
      | (~ alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp))) | FpCmp_8U_23U_true_if_acc_10_itm_8));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1 = (fsm_output[1]) & (~((~(FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1
      | (~ alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp))) | FpCmp_8U_23U_true_if_acc_8_itm_8));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2 = (fsm_output[1]) & (~((~(FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1
      | (~ alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp))) | FpCmp_8U_23U_true_if_acc_6_itm_8));
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3 = (fsm_output[1]) & (~((~(FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1
      | (~ alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp))) | FpCmp_8U_23U_true_if_acc_4_itm_8));
  assign alu_loop_op_else_else_if_and_cse = (fsm_output[1]) & ((cfg_alu_algo_1_sva_2!=2'b00));
  assign alu_loop_op_else_else_if_and_1_cse = (fsm_output[1]) & (cfg_alu_algo_1_sva_2[0]);
  assign FpAdd_8U_23U_if_2_and_tmp = (fsm_output[1]) & reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse;
  assign FpAdd_8U_23U_if_2_and_tmp_1 = (fsm_output[1]) & reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse;
  assign FpAdd_8U_23U_if_2_and_tmp_2 = (fsm_output[1]) & reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse;
  assign FpAdd_8U_23U_if_2_and_tmp_3 = (fsm_output[1]) & reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse;
  assign or_dcpl = (nor_397_cse & (~ FpAlu_8U_23U_equal_tmp_23) & FpAlu_8U_23U_nor_dfs_6)
      | io_read_cfg_alu_bypass_rsc_svs_8;
  assign mux_tmp = MUX_s_1_2_2(FpNormalize_8U_49U_oelse_not_9, alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1,
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]);
  assign mux_tmp_348 = MUX_s_1_2_2(FpNormalize_8U_49U_oelse_not_11, alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1,
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]);
  assign mux_tmp_349 = MUX_s_1_2_2(FpNormalize_8U_49U_oelse_not_13, alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1,
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]);
  assign mux_tmp_350 = MUX_s_1_2_2(FpNormalize_8U_49U_oelse_not_15, alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1,
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]);
  assign or_dcpl_272 = FpAlu_8U_23U_equal_tmp_29 | FpAlu_8U_23U_equal_tmp_26;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_iswt0 <= 1'b0;
      reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      chn_alu_out_rsci_iswt0 <= 1'b0;
      chn_alu_op_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_alu_in_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse <= or_tmp_695;
      chn_alu_out_rsci_iswt0 <= and_dcpl_43;
      chn_alu_op_rsci_iswt0 <= and_357_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_alu_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_alu_in_rsci_ld_core_psct <= chn_alu_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_0 <= 1'b0;
      chn_alu_out_rsci_d_32 <= 1'b0;
      chn_alu_out_rsci_d_96 <= 1'b0;
    end
    else if ( chn_alu_out_and_cse ) begin
      chn_alu_out_rsci_d_0 <= MUX_s_1_2_2((reg_AluIn_data_sva_4_30_0_1_itm[0]), (alu_loop_op_mux_209_nl),
          and_dcpl_40);
      chn_alu_out_rsci_d_32 <= MUX_s_1_2_2((reg_AluIn_data_sva_4_62_32_1_itm[0]),
          (alu_loop_op_mux_210_nl), and_dcpl_40);
      chn_alu_out_rsci_d_96 <= MUX_s_1_2_2((reg_AluIn_data_sva_4_126_96_1_itm[0]),
          (alu_loop_op_mux_212_nl), and_dcpl_40);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_22_1 <= 22'b0;
      chn_alu_out_rsci_d_54_33 <= 22'b0;
    end
    else if ( and_734_cse ) begin
      chn_alu_out_rsci_d_22_1 <= MUX1HOT_v_22_3_2((FpAlu_8U_23U_and_5_nl), AluOut_data_2_22_1_lpi_1_dfm_3,
          (reg_AluIn_data_sva_4_30_0_1_itm[22:1]), {nor_437_cse , asn_267 , or_dcpl});
      chn_alu_out_rsci_d_54_33 <= MUX1HOT_v_22_3_2((FpAlu_8U_23U_and_8_nl), IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4,
          (reg_AluIn_data_sva_4_62_32_1_itm[22:1]), {nor_437_cse , asn_267 , or_dcpl});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_30_23 <= 8'b0;
      chn_alu_out_rsci_d_31 <= 1'b0;
      chn_alu_out_rsci_d_62_55 <= 8'b0;
      chn_alu_out_rsci_d_63 <= 1'b0;
      chn_alu_out_rsci_d_95 <= 1'b0;
      chn_alu_out_rsci_d_118_97 <= 22'b0;
      chn_alu_out_rsci_d_126_119 <= 8'b0;
      chn_alu_out_rsci_d_127 <= 1'b0;
    end
    else if ( chn_alu_out_and_1_cse ) begin
      chn_alu_out_rsci_d_30_23 <= MUX1HOT_v_8_3_2((FpAlu_8U_23U_and_4_nl), AluOut_data_2_30_23_lpi_1_dfm_3,
          reg_AluIn_data_sva_4_30_0_itm, {(nor_406_nl) , asn_267 , or_996_tmp});
      chn_alu_out_rsci_d_31 <= mux_177_itm_4;
      chn_alu_out_rsci_d_62_55 <= MUX1HOT_v_8_3_2((FpAlu_8U_23U_and_7_nl), FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13,
          reg_AluIn_data_sva_4_62_32_itm, {(nor_407_nl) , asn_267 , or_997_tmp});
      chn_alu_out_rsci_d_63 <= mux_181_itm_4;
      chn_alu_out_rsci_d_95 <= AluOut_data_2_31_lpi_1_dfm_7;
      chn_alu_out_rsci_d_118_97 <= MUX1HOT_v_22_3_2(FpAlu_8U_23U_o_22_1_lpi_1_dfm_2,
          IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4, (reg_AluIn_data_sva_4_126_96_1_itm[22:1]),
          {nor_397_cse , asn_267 , io_read_cfg_alu_bypass_rsc_svs_8});
      chn_alu_out_rsci_d_126_119 <= MUX1HOT_v_8_3_2(FpAlu_8U_23U_o_30_23_lpi_1_dfm_2,
          FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13, reg_AluIn_data_sva_4_126_96_itm, {nor_397_cse
          , asn_267 , io_read_cfg_alu_bypass_rsc_svs_8});
      chn_alu_out_rsci_d_127 <= mux_189_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_64 <= 1'b0;
    end
    else if ( chn_alu_out_and_8_cse & chn_alu_out_or_cse ) begin
      chn_alu_out_rsci_d_64 <= MUX_s_1_2_2((reg_AluIn_data_sva_4_94_64_1_itm[0]),
          alu_loop_op_mux_204_mx1w1, and_dcpl_40);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_out_rsci_d_86_65 <= 22'b0;
      chn_alu_out_rsci_d_94_87 <= 8'b0;
    end
    else if ( chn_alu_out_and_18_cse ) begin
      chn_alu_out_rsci_d_86_65 <= AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0;
      chn_alu_out_rsci_d_94_87 <= AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_alu_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_43 | and_dcpl_45) ) begin
      reg_chn_alu_out_rsci_ld_core_psct_cse <= ~ and_dcpl_45;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_alu_op_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & (and_357_cse | (and_dcpl_30 & and_dcpl_46 & cfg_alu_src_1_sva_st_1
        & cfg_alu_src_rsci_d) | chn_alu_op_rsci_ld_core_psct_mx0c1) ) begin
      chn_alu_op_rsci_ld_core_psct <= ~ chn_alu_op_rsci_ld_core_psct_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_695 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluIn_data_sva_127 <= 128'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
      io_read_cfg_alu_bypass_rsc_svs_5 <= 1'b0;
    end
    else if ( AluIn_data_and_cse ) begin
      AluIn_data_sva_127 <= chn_alu_in_rsci_d_mxwt;
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0;
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0;
      io_read_cfg_alu_bypass_rsc_svs_5 <= cfg_alu_bypass_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_28 <= 2'b0;
    end
    else if ( core_wen & cfg_alu_algo_cfg_alu_algo_or_3_cse & (~ (mux_23_nl)) ) begin
      cfg_alu_algo_1_sva_st_28 <= cfg_alu_algo_cfg_alu_algo_mux_3_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_cfg_alu_algo_1_sva_st_13_cse <= 2'b0;
    end
    else if ( core_wen & cfg_alu_algo_cfg_alu_algo_or_3_cse & (~ (mux_31_nl)) ) begin
      reg_cfg_alu_algo_1_sva_st_13_cse <= cfg_alu_algo_cfg_alu_algo_mux_3_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_22 <= 2'b0;
    end
    else if ( core_wen & cfg_alu_algo_cfg_alu_algo_or_3_cse & (~ mux_34_itm) ) begin
      cfg_alu_algo_1_sva_st_22 <= MUX_v_2_2_2(cfg_alu_algo_rsci_d, cfg_alu_algo_1_sva_st,
          and_dcpl_81);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_op_1_sva_1 <= 32'b0;
    end
    else if ( chn_alu_out_and_8_cse & (and_dcpl_83 | and_167_rgt) & (mux_38_nl) )
        begin
      cfg_alu_op_1_sva_1 <= MUX_v_32_2_2(cfg_alu_op_rsci_d, (chn_alu_op_rsci_d_mxwt[127:96]),
          and_167_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_src_1_sva_st_1 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_83 & (fsm_output[1])) | (and_dcpl_30 & and_dcpl_46
        & cfg_alu_src_1_sva_st_1) | cfg_alu_src_1_sva_st_1_mx0c1) ) begin
      cfg_alu_src_1_sva_st_1 <= MUX_s_1_2_2(cfg_alu_src_rsci_d, cfg_alu_src_1_sva_st,
          cfg_alu_src_1_sva_st_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      io_read_cfg_alu_bypass_rsc_svs_st_1 <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_35 | and_dcpl_32 | (~ chn_alu_in_rsci_bawt)
        | (fsm_output[0]))) ) begin
      io_read_cfg_alu_bypass_rsc_svs_st_1 <= cfg_alu_bypass_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_64 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6 <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6 <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2;
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6 <= FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6 <= FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1;
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6 <= FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= IsNaN_8U_23U_4_nor_3_itm_3;
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1;
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6 <= FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= IsNaN_8U_23U_4_nor_2_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse
          <= 1'b0;
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5 <= 8'b0;
      reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5 <= 8'b0;
      reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5 <= 8'b0;
      reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse
          <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5 <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_8_cse ) begin
      reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse
          <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st,
          and_dcpl_99);
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm, and_dcpl_99);
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm, and_dcpl_99);
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm, and_dcpl_99);
      reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse
          <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st,
          and_dcpl_99);
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm, and_dcpl_99);
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm, and_dcpl_99);
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm, and_dcpl_99);
      reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse
          <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st,
          and_dcpl_99);
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm, and_dcpl_99);
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm, and_dcpl_99);
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm, and_dcpl_99);
      reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse
          <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st,
          and_dcpl_99);
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0,
          alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm, and_dcpl_99);
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm, and_dcpl_99);
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5 <= MUX_v_8_2_2(FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0,
          FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_3_lpi_1_dfm_2_30_0_1 <= 31'b0;
      else_AluOp_data_2_lpi_1_dfm_2_30_0_1 <= 31'b0;
      else_AluOp_data_1_lpi_1_dfm_2_30_0_1 <= 31'b0;
      else_AluOp_data_0_lpi_1_dfm_2_30_0_1 <= 31'b0;
      cfg_alu_algo_1_sva_st_23 <= 2'b0;
    end
    else if ( else_AluOp_data_and_10_cse ) begin
      else_AluOp_data_3_lpi_1_dfm_2_30_0_1 <= MUX_v_31_2_2((chn_alu_op_rsci_d_mxwt[126:96]),
          (cfg_alu_op_1_sva_1[30:0]), else_AluOp_data_else_AluOp_data_nor_nl);
      else_AluOp_data_2_lpi_1_dfm_2_30_0_1 <= else_AluOp_data_2_lpi_1_dfm_mx0[30:0];
      else_AluOp_data_1_lpi_1_dfm_2_30_0_1 <= else_AluOp_data_1_lpi_1_dfm_mx0[30:0];
      else_AluOp_data_0_lpi_1_dfm_2_30_0_1 <= else_AluOp_data_0_lpi_1_dfm_mx0[30:0];
      cfg_alu_algo_1_sva_st_23 <= cfg_alu_algo_1_sva_st_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluIn_data_sva_128 <= 128'b0;
      io_read_cfg_alu_bypass_rsc_svs_st_5 <= 1'b0;
      alu_loop_op_unequal_tmp_6 <= 1'b0;
      io_read_cfg_alu_bypass_rsc_svs_6 <= 1'b0;
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( AluIn_data_and_1_cse ) begin
      AluIn_data_sva_128 <= AluIn_data_sva_127;
      io_read_cfg_alu_bypass_rsc_svs_st_5 <= io_read_cfg_alu_bypass_rsc_svs_st_1;
      alu_loop_op_unequal_tmp_6 <= ~((cfg_precision==2'b10));
      io_read_cfg_alu_bypass_rsc_svs_6 <= io_read_cfg_alu_bypass_rsc_svs_5;
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_96 | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_7 <= 8'b0;
      FpAdd_8U_23U_qr_3_lpi_1_dfm_7 <= 8'b0;
      FpAdd_8U_23U_qr_4_lpi_1_dfm_7 <= 8'b0;
      FpAdd_8U_23U_qr_lpi_1_dfm_7 <= 8'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_and_39_cse ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_7 <= FpAdd_8U_23U_qr_2_lpi_1_dfm_6;
      FpAdd_8U_23U_qr_3_lpi_1_dfm_7 <= FpAdd_8U_23U_qr_3_lpi_1_dfm_6;
      FpAdd_8U_23U_qr_4_lpi_1_dfm_7 <= FpAdd_8U_23U_qr_4_lpi_1_dfm_6;
      FpAdd_8U_23U_qr_lpi_1_dfm_7 <= FpAdd_8U_23U_qr_lpi_1_dfm_6;
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_lpi_1_dfm_st_4;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5 <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5 <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5 <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5 <= 50'b0;
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2 <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_4_cse ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5 <= MUX_v_50_2_2(z_out_12, FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm,
          FpAdd_8U_23U_int_mant_p1_or_3_cse);
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5 <= MUX_v_50_2_2(z_out_13, FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm,
          FpAdd_8U_23U_int_mant_p1_or_3_cse);
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5 <= MUX_v_50_2_2(z_out_14, FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm,
          FpAdd_8U_23U_int_mant_p1_or_3_cse);
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5 <= MUX_v_50_2_2(z_out_15, FpAdd_8U_23U_int_mant_p1_lpi_1_dfm,
          FpAdd_8U_23U_int_mant_p1_or_3_cse);
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2 <= MUX_s_1_2_2((z_out_15[49]),
          alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm, and_dcpl_99);
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= MUX_s_1_2_2((z_out_14[49]),
          alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm, and_dcpl_99);
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2 <= MUX_s_1_2_2((z_out_13[49]),
          alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm, and_dcpl_99);
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= MUX_s_1_2_2((z_out_12[49]),
          alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_59_nl) ) begin
      FpNormalize_8U_49U_if_or_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_itm_mx0w0,
          FpNormalize_8U_49U_if_or_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_61_nl) ) begin
      FpNormalize_8U_49U_if_or_1_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_1_itm_mx0w0,
          FpNormalize_8U_49U_if_or_1_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_2_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_63_nl) ) begin
      FpNormalize_8U_49U_if_or_2_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_2_itm_mx0w0,
          FpNormalize_8U_49U_if_or_2_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_65_nl) ) begin
      FpNormalize_8U_49U_if_or_3_itm_2 <= MUX_s_1_2_2(FpNormalize_8U_49U_if_or_3_itm_mx0w0,
          FpNormalize_8U_49U_if_or_3_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_24 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_67_nl) ) begin
      cfg_alu_algo_1_sva_st_24 <= cfg_alu_algo_1_sva_st_23;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      io_read_cfg_alu_bypass_rsc_svs_st_6 <= 1'b0;
      AluIn_data_sva_3_62_32_1 <= 31'b0;
      AluIn_data_sva_3_30_0_1 <= 31'b0;
      AluIn_data_sva_3_94_64_1 <= 31'b0;
      AluIn_data_sva_3_126_96_1 <= 31'b0;
      alu_loop_op_unequal_tmp_7 <= 1'b0;
      io_read_cfg_alu_bypass_rsc_svs_7 <= 1'b0;
    end
    else if ( and_550_cse ) begin
      io_read_cfg_alu_bypass_rsc_svs_st_6 <= io_read_cfg_alu_bypass_rsc_svs_st_5;
      AluIn_data_sva_3_62_32_1 <= AluIn_data_sva_128[62:32];
      AluIn_data_sva_3_30_0_1 <= AluIn_data_sva_128[30:0];
      AluIn_data_sva_3_94_64_1 <= AluIn_data_sva_128[94:64];
      AluIn_data_sva_3_126_96_1 <= AluIn_data_sva_128[126:96];
      alu_loop_op_unequal_tmp_7 <= alu_loop_op_unequal_tmp_6;
      io_read_cfg_alu_bypass_rsc_svs_7 <= io_read_cfg_alu_bypass_rsc_svs_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & ((or_1087_cse & main_stage_v_3) | main_stage_v_4_mx0c1)
        ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 <= 8'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse & (mux_74_nl)
        ) begin
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 <= MUX_v_8_2_2(FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0,
          IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3, and_dcpl_108);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 <= 8'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse & (mux_80_nl)
        ) begin
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 <= MUX_v_8_2_2(FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0,
          IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3, and_dcpl_108);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 <= 8'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse & (mux_86_nl)
        ) begin
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 <= MUX_v_8_2_2(FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0,
          IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3, and_dcpl_108);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_lpi_1_dfm_13 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_92_nl) ) begin
      FpAdd_8U_23U_o_expo_lpi_1_dfm_13 <= FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_94_nl) ) begin
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3
          <= MUX_s_1_2_2(alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1, alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2,
          and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_96_nl) ) begin
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3
          <= MUX_s_1_2_2(alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1, alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2,
          and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_98_nl) ) begin
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3
          <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1, alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2,
          and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_100_nl) ) begin
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3
          <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1, alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2,
          and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_126_96_itm <= 8'b0;
    end
    else if ( ((nand_109_cse & FpAlu_8U_23U_nor_dfs_5 & nor_430_cse & IsNaN_8U_23U_land_lpi_1_dfm_10)
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_126_96_itm <= AluIn_data_mux1h_7_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_126_96_1_itm <= 23'b0;
    end
    else if ( (((and_564_cse | ((~ FpAlu_8U_23U_equal_tmp_22) & IsNaN_8U_23U_land_lpi_1_dfm_10))
        & FpAlu_8U_23U_nor_dfs_5 & (~ alu_loop_op_unequal_tmp_7) & (~ io_read_cfg_alu_bypass_rsc_svs_st_6))
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_126_96_1_itm <= AluIn_data_mux1h_7_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_8_cse ) begin
      IsNaN_8U_23U_land_lpi_1_dfm_11 <= IsNaN_8U_23U_land_lpi_1_dfm_10;
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 <= IsNaN_8U_23U_land_3_lpi_1_dfm_10;
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 <= IsNaN_8U_23U_land_2_lpi_1_dfm_10;
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 <= IsNaN_8U_23U_land_1_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= 1'b0;
      FpAdd_8U_23U_and_2_tmp_3 <= 1'b0;
      FpAdd_8U_23U_and_1_tmp_3 <= 1'b0;
      FpAdd_8U_23U_and_tmp_2 <= 1'b0;
      FpAdd_8U_23U_and_3_tmp_3 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_aelse_and_cse ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_lpi_1_dfm_8;
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
      FpAdd_8U_23U_and_2_tmp_3 <= alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1
          & alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
      FpAdd_8U_23U_and_1_tmp_3 <= alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1
          & alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
      FpAdd_8U_23U_and_tmp_2 <= alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
          & alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
      FpAdd_8U_23U_and_3_tmp_3 <= alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1
          & alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2 <= 1'b0;
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2 <= 1'b0;
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2 <= 1'b0;
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_else_and_4_cse ) begin
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2 <= MUX_s_1_2_2(alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp,
          alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st, and_dcpl_99);
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2 <= MUX_s_1_2_2(alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp,
          alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st, and_dcpl_99);
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2 <= MUX_s_1_2_2(alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp,
          alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st, and_dcpl_99);
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2 <= MUX_s_1_2_2(alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp,
          alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_94_64_itm <= 8'b0;
    end
    else if ( ((nand_109_cse & FpAlu_8U_23U_nor_dfs_5 & nor_430_cse & IsNaN_8U_23U_land_3_lpi_1_dfm_10)
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_94_64_itm <= AluIn_data_mux1h_9_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_94_64_1_itm <= 23'b0;
    end
    else if ( (((and_564_cse | ((~ FpAlu_8U_23U_equal_tmp_22) & IsNaN_8U_23U_land_3_lpi_1_dfm_10))
        & FpAlu_8U_23U_nor_dfs_5 & (~ alu_loop_op_unequal_tmp_7) & (~ io_read_cfg_alu_bypass_rsc_svs_st_6))
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_94_64_1_itm <= AluIn_data_mux1h_9_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_62_32_itm <= 8'b0;
    end
    else if ( ((nand_109_cse & FpAlu_8U_23U_nor_dfs_5 & nor_430_cse & IsNaN_8U_23U_land_2_lpi_1_dfm_10)
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_62_32_itm <= AluIn_data_mux1h_11_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_62_32_1_itm <= 23'b0;
    end
    else if ( (((and_564_cse | ((~ FpAlu_8U_23U_equal_tmp_22) & IsNaN_8U_23U_land_2_lpi_1_dfm_10))
        & FpAlu_8U_23U_nor_dfs_5 & (~ alu_loop_op_unequal_tmp_7) & (~ io_read_cfg_alu_bypass_rsc_svs_st_6))
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_62_32_1_itm <= AluIn_data_mux1h_11_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_30_0_itm <= 8'b0;
    end
    else if ( ((nand_109_cse & FpAlu_8U_23U_nor_dfs_5 & nor_430_cse & IsNaN_8U_23U_land_1_lpi_1_dfm_10)
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_30_0_itm <= AluIn_data_mux1h_13_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_AluIn_data_sva_4_30_0_1_itm <= 23'b0;
    end
    else if ( (((and_564_cse | ((~ FpAlu_8U_23U_equal_tmp_22) & IsNaN_8U_23U_land_1_lpi_1_dfm_10))
        & FpAlu_8U_23U_nor_dfs_5 & (~ alu_loop_op_unequal_tmp_7) & (~ io_read_cfg_alu_bypass_rsc_svs_st_6))
        | io_read_cfg_alu_bypass_rsc_svs_7) & and_dcpl & or_1087_cse ) begin
      reg_AluIn_data_sva_4_30_0_1_itm <= AluIn_data_mux1h_13_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_nor_dfs_6 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_26 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_23 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_29 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_32 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_82_cse ) begin
      FpAlu_8U_23U_nor_dfs_6 <= FpAlu_8U_23U_nor_dfs_5;
      FpAlu_8U_23U_equal_tmp_26 <= FpAlu_8U_23U_equal_tmp_25;
      FpAlu_8U_23U_equal_tmp_23 <= FpAlu_8U_23U_equal_tmp_22;
      FpAlu_8U_23U_equal_tmp_29 <= FpAlu_8U_23U_equal_tmp_28;
      FpAlu_8U_23U_equal_tmp_32 <= FpAlu_8U_23U_equal_tmp_31;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1 <= 31'b0;
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1 <= 31'b0;
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1 <= 31'b0;
    end
    else if ( FpCmp_8U_23U_true_o_and_cse ) begin
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1 <= FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1;
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1 <= FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1;
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1 <= FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_22_1_lpi_1_dfm_3 <= 22'b0;
    end
    else if ( ((((mux_383_nl) | io_read_cfg_alu_bypass_rsc_svs_8) & main_stage_v_4)
        | nor_tmp_144) & or_1087_cse & core_wen ) begin
      AluOut_data_2_22_1_lpi_1_dfm_3 <= MUX_v_22_2_2(AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0,
          IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2, and_dcpl_127);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_127_nl)) ) begin
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1 <= FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_1087_cse & alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp)
        | and_211_rgt) & (~ mux_109_itm) ) begin
      FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8 <= MUX_s_1_2_2(FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0,
          nor_41_cse, and_211_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_128_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_30_23_lpi_1_dfm_3 <= 8'b0;
    end
    else if ( (((FpAlu_8U_23U_equal_tmp_29 | FpAlu_8U_23U_equal_tmp_26 | FpAlu_8U_23U_nor_dfs_6
        | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8)
        & main_stage_v_4) | nor_tmp_144) & or_1087_cse & core_wen ) begin
      AluOut_data_2_30_23_lpi_1_dfm_3 <= MUX_v_8_2_2(AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0,
          IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2, and_dcpl_127);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1 <= 31'b0;
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1 <= 31'b0;
    end
    else if ( FpCmp_8U_23U_false_o_and_1_cse ) begin
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1 <= FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1;
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1 <= FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_1087_cse & alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp)
        | and_213_rgt) & (~ mux_109_itm) ) begin
      FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8 <= MUX_s_1_2_2(FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0,
          nor_37_cse, and_213_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_130_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_1087_cse & alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp)
        | and_215_rgt) & (~ mux_109_itm) ) begin
      FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8 <= MUX_s_1_2_2(FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0,
          nor_33_cse, and_215_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_131_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_133_nl)) ) begin
      FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1 <= FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_0_sva_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_135_nl)) ) begin
      FpAlu_8U_23U_o_0_sva_9 <= FpAlu_8U_23U_o_0_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_0_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( (~((~(FpAlu_8U_23U_equal_tmp_29 | FpAlu_8U_23U_equal_tmp_23 | FpAlu_8U_23U_equal_tmp_26
        | FpAlu_8U_23U_nor_dfs_6)) | alu_loop_op_unequal_tmp_8)) & (~ io_read_cfg_alu_bypass_rsc_svs_8)
        & main_stage_v_4 & core_wen & or_1087_cse ) begin
      FpAlu_8U_23U_o_0_lpi_1_dfm_4 <= FpAlu_8U_23U_o_0_lpi_1_dfm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_136_nl)) ) begin
      FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1 <= FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_22_1_lpi_1_dfm_4 <= 22'b0;
      FpAlu_8U_23U_o_30_23_lpi_1_dfm_4 <= 8'b0;
    end
    else if ( and_524_cse ) begin
      FpAlu_8U_23U_o_22_1_lpi_1_dfm_4 <= FpAlu_8U_23U_o_22_1_lpi_1_dfm_2;
      FpAlu_8U_23U_o_30_23_lpi_1_dfm_4 <= FpAlu_8U_23U_o_30_23_lpi_1_dfm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_inf_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_1087_cse & alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp)
        | and_217_rgt) & (~ mux_109_itm) ) begin
      FpAdd_8U_23U_is_inf_lpi_1_dfm_8 <= MUX_s_1_2_2(FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0,
          nor_45_cse, and_217_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3 <= 8'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_137_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_35 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_138_nl)) ) begin
      FpAlu_8U_23U_equal_tmp_35 <= FpAlu_8U_23U_equal_tmp_34;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_25 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_139_nl)) ) begin
      cfg_alu_algo_1_sva_st_25 <= cfg_alu_algo_1_sva_st_24;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      mux_189_itm_4 <= 1'b0;
      alu_loop_op_unequal_tmp_8 <= 1'b0;
      io_read_cfg_alu_bypass_rsc_svs_8 <= 1'b0;
      mux_177_itm_4 <= 1'b0;
      AluOut_data_2_31_lpi_1_dfm_7 <= 1'b0;
      mux_181_itm_4 <= 1'b0;
      io_read_cfg_alu_bypass_rsc_svs_st_7 <= 1'b0;
    end
    else if ( and_cse ) begin
      mux_189_itm_4 <= mux_189_itm_3;
      alu_loop_op_unequal_tmp_8 <= alu_loop_op_unequal_tmp_7;
      io_read_cfg_alu_bypass_rsc_svs_8 <= io_read_cfg_alu_bypass_rsc_svs_7;
      mux_177_itm_4 <= mux_177_itm_3;
      AluOut_data_2_31_lpi_1_dfm_7 <= AluOut_data_2_31_lpi_1_dfm_6;
      mux_181_itm_4 <= mux_181_itm_3;
      io_read_cfg_alu_bypass_rsc_svs_st_7 <= io_read_cfg_alu_bypass_rsc_svs_st_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_0_0_sva_11 <= 1'b0;
      AluOut_data_1_0_sva_12 <= 1'b0;
    end
    else if ( AluOut_data_and_8_cse ) begin
      AluOut_data_0_0_sva_11 <= AluOut_data_0_0_sva_10;
      AluOut_data_1_0_sva_12 <= AluOut_data_1_0_sva_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4 <= 22'b0;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4 <= 22'b0;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4 <= 22'b0;
    end
    else if ( IntSaturation_33U_32U_and_cse ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4 <= IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_0_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( (mux_362_nl) & core_wen ) begin
      AluOut_data_2_0_lpi_1_dfm_3 <= MUX1HOT_s_1_3_2((reg_AluIn_data_sva_4_94_64_1_itm[0]),
          alu_loop_op_mux_204_mx1w1, AluOut_data_2_0_sva_10, {(and_218_nl) , (and_220_nl)
          , and_dcpl_127});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_0_sva_11 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse & (~ mux_143_itm)
        ) begin
      AluOut_data_2_0_sva_11 <= MUX_s_1_2_2(AluOut_data_2_0_sva_10, FpAlu_8U_23U_o_0_sva_8,
          and_dcpl_108);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_85) & (mux_145_nl) ) begin
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2
          <= alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_85) & (mux_146_nl) ) begin
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2
          <= alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_85) & (mux_147_nl) ) begin
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2
          <= alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_85) & (mux_148_nl) ) begin
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2
          <= alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st <= 1'b0;
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st <= 1'b0;
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st <= 1'b0;
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_else_and_cse ) begin
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st <= alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st <= alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st <= alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st <= alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_150_nl) ) begin
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_152_nl) ) begin
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_154_nl) ) begin
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_156_nl) ) begin
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= IsNaN_8U_23U_1_land_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_itm <= 1'b0;
    end
    else if ( chn_alu_out_and_8_cse & (~ or_dcpl_89) & (mux_157_nl) ) begin
      FpNormalize_8U_49U_if_or_itm <= FpNormalize_8U_49U_if_or_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm <= 50'b0;
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm <= 50'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_12_cse ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm <= z_out_12;
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm <= z_out_13;
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm <= z_out_14;
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm <= z_out_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_1_itm <= 1'b0;
    end
    else if ( chn_alu_out_and_8_cse & (~ or_dcpl_89) & (mux_158_nl) ) begin
      FpNormalize_8U_49U_if_or_1_itm <= FpNormalize_8U_49U_if_or_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_2_itm <= 1'b0;
    end
    else if ( chn_alu_out_and_8_cse & (~ or_dcpl_89) & (mux_159_nl) ) begin
      FpNormalize_8U_49U_if_or_2_itm <= FpNormalize_8U_49U_if_or_2_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_8U_49U_if_or_3_itm <= 1'b0;
    end
    else if ( chn_alu_out_and_8_cse & (~ or_dcpl_89) & (mux_160_nl) ) begin
      FpNormalize_8U_49U_if_or_3_itm <= FpNormalize_8U_49U_if_or_3_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
    end
    else if ( FpAdd_8U_23U_if_3_and_cse ) begin
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm <= z_out_15[49];
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= z_out_14[49];
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm <= z_out_13[49];
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= z_out_12[49];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
    end
    else if ( IsZero_8U_23U_and_4_cse ) begin
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= MUX_s_1_2_2(alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3, and_dcpl_81);
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= MUX_s_1_2_2(alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0,
          alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3, and_dcpl_81);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm <= 8'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm <= 8'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm <= 8'b0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm <= 8'b0;
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm <= 8'b0;
    end
    else if ( IsZero_8U_23U_1_and_cse ) begin
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm <= FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0;
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm <= FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm <= FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0;
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm <= FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm <= FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0;
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm <= FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0;
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm <= FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0;
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm <= FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st
          <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st
          <= 1'b0;
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_cse ) begin
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st
          <= alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st
          <= alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st
          <= alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0;
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st
          <= alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st_20 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_109) & (~ (mux_172_nl)) ) begin
      cfg_alu_algo_1_sva_st_20 <= cfg_alu_algo_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_st <= 2'b0;
    end
    else if ( core_wen & (~(or_dcpl_109 | (fsm_output[0]))) ) begin
      cfg_alu_algo_1_sva_st <= cfg_alu_algo_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_src_1_sva_st <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_35 | or_tmp_386 | and_dcpl_32 | (fsm_output[0])))
        ) begin
      cfg_alu_src_1_sva_st <= cfg_alu_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_alu_algo_1_sva_2 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_49) & (~ mux_34_itm) ) begin
      cfg_alu_algo_1_sva_2 <= cfg_alu_algo_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_6 <= 8'b0;
    end
    else if ( core_wen & (and_231_rgt | and_233_rgt | and_dcpl_99) & not_tmp_29 )
        begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm_6 <= MUX1HOT_v_8_3_2((AluIn_data_sva_127[30:23]),
          else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23, FpAdd_8U_23U_qr_2_lpi_1_dfm,
          {and_231_rgt , and_233_rgt , and_dcpl_99});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_6 <= 8'b0;
    end
    else if ( core_wen & (and_235_rgt | and_237_rgt | and_dcpl_99) & not_tmp_29 )
        begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm_6 <= MUX1HOT_v_8_3_2((AluIn_data_sva_127[62:55]),
          else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23, FpAdd_8U_23U_qr_3_lpi_1_dfm,
          {and_235_rgt , and_237_rgt , and_dcpl_99});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_6 <= 8'b0;
    end
    else if ( core_wen & (and_239_rgt | and_241_rgt | and_dcpl_99) & not_tmp_29 )
        begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm_6 <= MUX1HOT_v_8_3_2((AluIn_data_sva_127[94:87]),
          else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23, FpAdd_8U_23U_qr_4_lpi_1_dfm,
          {and_239_rgt , and_241_rgt , and_dcpl_99});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm_6 <= 8'b0;
    end
    else if ( core_wen & (and_243_rgt | and_245_rgt | and_dcpl_99) & not_tmp_29 )
        begin
      FpAdd_8U_23U_qr_lpi_1_dfm_6 <= MUX1HOT_v_8_3_2((AluIn_data_sva_127[126:119]),
          else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23, FpAdd_8U_23U_qr_lpi_1_dfm, {and_243_rgt
          , and_245_rgt , and_dcpl_99});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_12_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= IsNaN_8U_23U_land_2_lpi_1_dfm_9;
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= IsNaN_8U_23U_land_1_lpi_1_dfm_9;
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= IsNaN_8U_23U_land_3_lpi_1_dfm_9;
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= IsNaN_8U_23U_land_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_0_sva_8 <= 1'b0;
    end
    else if ( core_wen & FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse & (~ (mux_182_nl))
        ) begin
      FpAlu_8U_23U_o_0_sva_8 <= MUX_s_1_2_2(FpAlu_8U_23U_o_0_sva_7, (IntSaturation_33U_32U_IntSaturation_33U_32U_or_nl),
          and_dcpl_165);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_0_sva_10 <= 1'b0;
      AluOut_data_1_0_sva_11 <= 1'b0;
      AluOut_data_0_0_sva_10 <= 1'b0;
    end
    else if ( AluOut_data_and_12_cse ) begin
      AluOut_data_2_0_sva_10 <= MUX_s_1_2_2(AluOut_data_2_0_sva_9, (IntSaturation_33U_32U_IntSaturation_33U_32U_or_3_nl),
          and_dcpl_165);
      AluOut_data_1_0_sva_11 <= MUX_s_1_2_2(AluOut_data_1_0_sva_10, (IntSaturation_33U_32U_IntSaturation_33U_32U_or_2_nl),
          and_dcpl_165);
      AluOut_data_0_0_sva_10 <= MUX_s_1_2_2(AluOut_data_0_0_sva_9, (IntSaturation_33U_32U_IntSaturation_33U_32U_or_1_nl),
          and_dcpl_165);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_22 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_25 <= 1'b0;
      FpAlu_8U_23U_nor_dfs_5 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_28 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_31 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_88_cse ) begin
      FpAlu_8U_23U_equal_tmp_22 <= FpAlu_8U_23U_equal_tmp_21;
      FpAlu_8U_23U_equal_tmp_25 <= FpAlu_8U_23U_equal_tmp_24;
      FpAlu_8U_23U_nor_dfs_5 <= FpAlu_8U_23U_nor_dfs_4;
      FpAlu_8U_23U_equal_tmp_28 <= FpAlu_8U_23U_equal_tmp_27;
      FpAlu_8U_23U_equal_tmp_31 <= FpAlu_8U_23U_equal_tmp_30;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_190_nl)) ) begin
      FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1 <= FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1 <= 31'b0;
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1 <= 31'b0;
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1 <= 31'b0;
    end
    else if ( FpCmp_8U_23U_true_o_and_5_cse ) begin
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1 <= FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1;
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1 <= FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1;
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1 <= FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_194_nl)) ) begin
      FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1 <= reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ (mux_196_nl)) ) begin
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1 <= reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1 <= 31'b0;
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1 <= 31'b0;
    end
    else if ( FpCmp_8U_23U_false_o_and_6_cse ) begin
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1 <= reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm;
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1 <= reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_34 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (~ mux_tmp_173) ) begin
      FpAlu_8U_23U_equal_tmp_34 <= FpAlu_8U_23U_equal_tmp_33;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3 <= 8'b0;
    end
    else if ( core_wen & IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse & (mux_200_nl)
        ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3 <= MUX1HOT_v_8_3_2((IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1[29:22]),
          (else_AluOp_data_2_lpi_1_dfm_2_30_0_1[30:23]), else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm,
          {and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3 <= 22'b0;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3 <= 22'b0;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3 <= 22'b0;
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2 <= 22'b0;
    end
    else if ( IntSaturation_33U_32U_and_11_cse ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3 <= IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1[21:0];
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3 <= IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1[21:0];
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3 <= IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1[21:0];
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2 <= IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1[21:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3 <= 8'b0;
    end
    else if ( core_wen & IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse & (mux_204_nl)
        ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3 <= MUX1HOT_v_8_3_2((IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1[29:22]),
          (else_AluOp_data_3_lpi_1_dfm_2_30_0_1[30:23]), else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm,
          {and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3 <= 8'b0;
    end
    else if ( core_wen & IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse & (mux_206_nl)
        ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3 <= MUX1HOT_v_8_3_2((IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1[29:22]),
          (else_AluOp_data_1_lpi_1_dfm_2_30_0_1[30:23]), else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm,
          {and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2 <= 8'b0;
    end
    else if ( core_wen & IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse & (mux_208_nl)
        ) begin
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2 <= MUX1HOT_v_8_3_2((IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1[29:22]),
          (else_AluOp_data_0_lpi_1_dfm_2_30_0_1[30:23]), else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm,
          {and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_31_lpi_1_dfm_6 <= 1'b0;
      mux_189_itm_3 <= 1'b0;
      mux_181_itm_3 <= 1'b0;
      mux_177_itm_3 <= 1'b0;
    end
    else if ( AluOut_data_and_15_cse ) begin
      AluOut_data_2_31_lpi_1_dfm_6 <= MUX1HOT_s_1_3_2((AluIn_data_sva_128[95]), (FpAlu_8U_23U_and_9_nl),
          (IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1[30]), {and_dcpl_170 , alu_loop_bypass_if_and_6_cse
          , alu_loop_bypass_if_and_7_cse});
      mux_189_itm_3 <= MUX1HOT_s_1_3_2((AluIn_data_sva_128[127]), (FpAlu_8U_23U_and_nl),
          (IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1[30]), {and_dcpl_170 , alu_loop_bypass_if_and_6_cse
          , alu_loop_bypass_if_and_7_cse});
      mux_181_itm_3 <= MUX1HOT_s_1_3_2((AluIn_data_sva_128[63]), FpAlu_8U_23U_and_6_itm_2,
          (IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1[30]), {and_dcpl_170 , alu_loop_bypass_if_and_6_cse
          , alu_loop_bypass_if_and_7_cse});
      mux_177_itm_3 <= MUX1HOT_s_1_3_2((AluIn_data_sva_128[31]), FpAlu_8U_23U_and_3_itm_2,
          (IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1[30]), {and_dcpl_170 , alu_loop_bypass_if_and_6_cse
          , alu_loop_bypass_if_and_7_cse});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_209_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2 <= MUX_v_23_2_2((else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0]),
          else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_210_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2 <= MUX_v_23_2_2((else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0]),
          else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_211_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2 <= MUX_v_23_2_2((else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0]),
          else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2 <= 23'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse
        & (mux_212_nl) ) begin
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2 <= MUX_v_23_2_2((else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0]),
          else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm, and_dcpl_99);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm <= 23'b0;
    end
    else if ( core_wen & (~(or_dcpl_127 | or_dcpl_125 | (cfg_alu_algo_1_sva_st_23[0])
        | IsNaN_8U_23U_land_1_lpi_1_dfm_st_4)) ) begin
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm <= else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm <= 23'b0;
    end
    else if ( core_wen & (~(or_dcpl_127 | or_dcpl_125 | (cfg_alu_algo_1_sva_st_23[0])
        | IsNaN_8U_23U_land_2_lpi_1_dfm_st_4)) ) begin
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm <= else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm <= 23'b0;
    end
    else if ( core_wen & (~(or_dcpl_127 | or_dcpl_125 | (cfg_alu_algo_1_sva_st_23[0])
        | IsNaN_8U_23U_land_3_lpi_1_dfm_st_4)) ) begin
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm <= else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm <= 23'b0;
    end
    else if ( core_wen & (~(or_dcpl_127 | or_dcpl_125 | (cfg_alu_algo_1_sva_st_23[0])
        | IsNaN_8U_23U_land_lpi_1_dfm_st_4)) ) begin
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm <= else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm <= 8'b0;
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm <= 8'b0;
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm <= 8'b0;
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm <= 8'b0;
    end
    else if ( FpAdd_8U_23U_int_mant_p1_and_cse ) begin
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm <= else_AluOp_data_2_lpi_1_dfm_2_30_0_1[30:23];
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm <= else_AluOp_data_1_lpi_1_dfm_2_30_0_1[30:23];
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm <= else_AluOp_data_0_lpi_1_dfm_2_30_0_1[30:23];
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm <= else_AluOp_data_3_lpi_1_dfm_2_30_0_1[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_21 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_24 <= 1'b0;
      FpAlu_8U_23U_nor_dfs_4 <= 1'b0;
      FpAlu_8U_23U_equal_tmp_27 <= 1'b0;
      FpAlu_8U_23U_and_3_itm_2 <= 1'b0;
      FpAlu_8U_23U_and_6_itm_2 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_94_cse ) begin
      FpAlu_8U_23U_equal_tmp_21 <= FpAlu_8U_23U_equal_tmp_1_mx0w0;
      FpAlu_8U_23U_equal_tmp_24 <= FpAlu_8U_23U_equal_tmp_mx0w0;
      FpAlu_8U_23U_nor_dfs_4 <= FpAlu_8U_23U_nor_dfs_mx0w0;
      FpAlu_8U_23U_equal_tmp_27 <= FpAlu_8U_23U_equal_tmp_2_mx0w0;
      FpAlu_8U_23U_and_3_itm_2 <= (FpAlu_8U_23U_mux1h_144_nl) & (~ FpAlu_8U_23U_equal_tmp_1_mx0w0);
      FpAlu_8U_23U_and_6_itm_2 <= (FpAlu_8U_23U_mux1h_148_nl) & (~ FpAlu_8U_23U_equal_tmp_1_mx0w0);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm <= 8'b0;
    end
    else if ( core_wen & ((and_dcpl_179 & and_dcpl_175 & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0
        & main_stage_v_1) | FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1) ) begin
      FpAdd_8U_23U_qr_2_lpi_1_dfm <= MUX_v_8_2_2((AluIn_data_sva_127[30:23]), else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23,
          FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm <= 8'b0;
    end
    else if ( core_wen & ((and_dcpl_179 & and_dcpl_175 & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0
        & main_stage_v_1) | FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1) ) begin
      FpAdd_8U_23U_qr_3_lpi_1_dfm <= MUX_v_8_2_2((AluIn_data_sva_127[62:55]), else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23,
          FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm <= 8'b0;
    end
    else if ( core_wen & ((and_dcpl_179 & and_dcpl_175 & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0
        & main_stage_v_1) | FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1) ) begin
      FpAdd_8U_23U_qr_4_lpi_1_dfm <= MUX_v_8_2_2((AluIn_data_sva_127[94:87]), else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23,
          FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm <= 8'b0;
    end
    else if ( core_wen & ((and_dcpl_179 & and_dcpl_175 & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0
        & main_stage_v_1) | FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1) ) begin
      FpAdd_8U_23U_qr_lpi_1_dfm <= MUX_v_8_2_2((AluIn_data_sva_127[126:119]), else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23,
          FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
    end
    else if ( IsZero_8U_23U_and_6_cse ) begin
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_16_cse ) begin
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= IsNaN_8U_23U_land_2_lpi_1_dfm_8;
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= IsNaN_8U_23U_land_1_lpi_1_dfm_8;
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= IsNaN_8U_23U_land_3_lpi_1_dfm_8;
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= IsNaN_8U_23U_land_lpi_1_dfm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_o_0_sva_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_218_nl) ) begin
      FpAlu_8U_23U_o_0_sva_7 <= FpAlu_8U_23U_o_0_sva_2_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_2_0_sva_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_219_nl) ) begin
      AluOut_data_2_0_sva_9 <= AluOut_data_2_0_sva_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      AluOut_data_1_0_sva_10 <= 1'b0;
      AluOut_data_0_0_sva_9 <= 1'b0;
    end
    else if ( AluOut_data_and_17_cse ) begin
      AluOut_data_1_0_sva_10 <= MUX1HOT_s_1_3_2(((AluIn_data_sva_127[63:32]) != else_AluOp_data_1_lpi_1_dfm_mx0),
          (alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0[0]), (alu_loop_op_else_else_else_else_ac_int_cctor_2_sva[0]),
          {(AluOut_data_or_1_nl) , (AluOut_data_or_2_nl) , (AluOut_data_and_7_nl)});
      AluOut_data_0_0_sva_9 <= MUX1HOT_s_1_3_2(((AluIn_data_sva_127[31:0]) != else_AluOp_data_0_lpi_1_dfm_mx0),
          (alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0[0]), (alu_loop_op_else_else_else_else_ac_int_cctor_1_sva[0]),
          {(AluOut_data_or_nl) , (AluOut_data_or_3_nl) , (AluOut_data_and_3_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_223_nl) ) begin
      FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1 <= FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1 <= 31'b0;
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1 <= 31'b0;
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1 <= 31'b0;
    end
    else if ( FpCmp_8U_23U_true_o_and_9_cse ) begin
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1 <= FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0[30:0];
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1 <= FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0[30:0];
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1 <= FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_30 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_225_nl) ) begin
      FpAlu_8U_23U_equal_tmp_30 <= FpAlu_8U_23U_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_equal_tmp_33 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_32) & (mux_226_nl) ) begin
      FpAlu_8U_23U_equal_tmp_33 <= FpAlu_8U_23U_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm <= 1'b0;
    end
    else if ( or_963_cse & core_wen & (~ alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2)
        & (~ io_read_cfg_alu_bypass_rsc_svs_5) & cfg_alu_algo_rsc_triosy_obj_bawt
        & or_1050_cse & and_dcpl_349 & cfg_alu_bypass_rsc_triosy_obj_bawt & (~ io_read_cfg_alu_bypass_rsc_svs_st_1)
        & or_1087_cse & main_stage_v_1 ) begin
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm <= alu_loop_op_else_o_mux1h_1_itm[31];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm <= 31'b0;
    end
    else if ( (~((mux_363_nl) | nor_202_cse)) & core_wen & (~ io_read_cfg_alu_bypass_rsc_svs_5)
        & and_dcpl_2 & and_dcpl_3 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1
        & or_1087_cse ) begin
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm <= alu_loop_op_else_o_mux1h_1_itm[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm <= 1'b0;
    end
    else if ( or_963_cse & core_wen & (~ alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2)
        & (~ io_read_cfg_alu_bypass_rsc_svs_5) & cfg_alu_algo_rsc_triosy_obj_bawt
        & or_1050_cse & and_dcpl_349 & cfg_alu_bypass_rsc_triosy_obj_bawt & (~ io_read_cfg_alu_bypass_rsc_svs_st_1)
        & or_1087_cse & main_stage_v_1 ) begin
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm <= alu_loop_op_else_o_mux1h_3_itm[31];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm <= 31'b0;
    end
    else if ( (~((mux_364_nl) | nor_202_cse)) & core_wen & (~ io_read_cfg_alu_bypass_rsc_svs_5)
        & and_dcpl_2 & and_dcpl_3 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1
        & or_1087_cse ) begin
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm <= alu_loop_op_else_o_mux1h_3_itm[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3
          <= 1'b0;
    end
    else if ( core_wen & ((or_1087_cse & (~ io_read_cfg_alu_bypass_rsc_svs_st_1))
        | and_293_rgt) & not_tmp_232 ) begin
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3
          <= MUX_s_1_2_2(alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2,
          and_293_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm <= 1'b0;
    end
    else if ( or_963_cse & core_wen & (~ alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2)
        & (~ io_read_cfg_alu_bypass_rsc_svs_5) & cfg_alu_algo_rsc_triosy_obj_bawt
        & or_1050_cse & and_dcpl_349 & cfg_alu_bypass_rsc_triosy_obj_bawt & (~ io_read_cfg_alu_bypass_rsc_svs_st_1)
        & or_1087_cse & main_stage_v_1 ) begin
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm <= alu_loop_op_else_o_mux1h_5_itm[31];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm <= 31'b0;
    end
    else if ( (~ (mux_365_nl)) & or_963_cse & core_wen & (~ io_read_cfg_alu_bypass_rsc_svs_5)
        & cfg_alu_algo_rsc_triosy_obj_bawt & cfg_alu_op_rsc_triosy_obj_bawt & and_dcpl_3
        & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1 & or_1087_cse
        ) begin
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm <= alu_loop_op_else_o_mux1h_5_itm[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm <= 1'b0;
    end
    else if ( core_wen & (~ io_read_cfg_alu_bypass_rsc_svs_5) & or_963_cse & and_dcpl_2
        & or_1050_cse & and_dcpl_3 & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1
        & (~(nor_269_cse | alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2)) )
        begin
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm <= alu_loop_op_else_o_mux1h_7_itm[31];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm <= 31'b0;
    end
    else if ( (~((mux_366_nl) | nor_202_cse)) & core_wen & (~ io_read_cfg_alu_bypass_rsc_svs_5)
        & cfg_alu_algo_rsc_triosy_obj_bawt & and_dcpl_349 & cfg_alu_bypass_rsc_triosy_obj_bawt
        & (~ io_read_cfg_alu_bypass_rsc_svs_st_1) & main_stage_v_1 & or_1087_cse
        ) begin
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm <= alu_loop_op_else_o_mux1h_7_itm[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2
          <= 1'b0;
      alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2
          <= 1'b0;
      alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2
          <= 1'b0;
    end
    else if ( IntSaturation_33U_32U_if_and_9_cse ) begin
      alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2
          <= alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2;
      alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2
          <= alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2;
      alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2
          <= alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAlu_8U_23U_mux1h_33_itm_2 <= 1'b0;
      FpAlu_8U_23U_mux1h_152_itm_2 <= 1'b0;
    end
    else if ( FpAlu_8U_23U_and_102_cse ) begin
      FpAlu_8U_23U_mux1h_33_itm_2 <= MUX1HOT_s_1_7_2((else_AluOp_data_3_lpi_1_dfm_mx0[31]),
          (AluIn_data_sva_127[127]), (FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0[31]), (FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0[31]),
          (alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0[0]), FpAlu_8U_23U_o_0_sva_2_mx0w0,
          (alu_loop_op_else_else_else_else_ac_int_cctor_sva[0]), {(FpAlu_8U_23U_and_74_nl)
          , (FpAlu_8U_23U_and_75_nl) , (FpAlu_8U_23U_and_76_nl) , (FpAlu_8U_23U_and_77_nl)
          , FpAlu_8U_23U_or_cse , (FpAlu_8U_23U_and_80_nl) , (FpAlu_8U_23U_and_81_nl)});
      FpAlu_8U_23U_mux1h_152_itm_2 <= MUX1HOT_s_1_7_2((else_AluOp_data_2_lpi_1_dfm_mx0[31]),
          (AluIn_data_sva_127[95]), (FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0[31]),
          (FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0[31]), (alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0[0]),
          AluOut_data_2_0_sva_3_mx0w0, (alu_loop_op_else_else_else_else_ac_int_cctor_3_sva[0]),
          {(FpAlu_8U_23U_and_66_nl) , (FpAlu_8U_23U_and_67_nl) , (FpAlu_8U_23U_and_68_nl)
          , (FpAlu_8U_23U_and_69_nl) , FpAlu_8U_23U_or_cse , (FpAlu_8U_23U_and_72_nl)
          , (FpAlu_8U_23U_and_73_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2
          <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_49) & (~ (mux_175_nl)) ) begin
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2
          <= cfg_alu_src_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2 <= 1'b0;
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_and_6_cse ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0, {and_dcpl_219 , and_dcpl_81
          , and_dcpl_222 , and_dcpl_225});
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0, {and_dcpl_219 , and_dcpl_81
          , and_dcpl_222 , and_dcpl_225});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 <= 1'b0;
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_and_cse ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm, IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0, {and_dcpl_219 , and_dcpl_81
          , and_dcpl_222 , and_dcpl_225});
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm, IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0, {and_dcpl_219 , and_dcpl_81
          , and_dcpl_222 , and_dcpl_225});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_20 | or_dcpl_46 | (cfg_alu_algo_1_sva_st_22!=2'b01)
        | and_dcpl_33 | io_read_cfg_alu_bypass_rsc_svs_st_1 | (~ main_stage_v_1)
        | or_dcpl_154)) & (~ (mux_277_nl)) ) begin
      FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2 <= FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_nor_3_itm_3 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse & (~ (mux_290_nl))
        ) begin
      IsNaN_8U_23U_4_nor_3_itm_3 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_2_nor_3_mx0w0, IsNaN_8U_23U_4_nor_3_itm_2,
          alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0, alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3,
          {and_dcpl_222 , and_dcpl_227 , and_dcpl_229 , and_dcpl_231});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_nor_2_itm_2 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse & (~ (mux_303_nl))
        ) begin
      IsNaN_8U_23U_4_nor_2_itm_2 <= MUX1HOT_s_1_4_2(IsNaN_8U_23U_2_nor_2_mx0w0, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm,
          alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2, IsNaN_8U_23U_4_nor_3_itm_2,
          {and_dcpl_222 , and_dcpl_227 , and_dcpl_229 , and_dcpl_231});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm <= 1'b0;
    end
    else if ( chn_alu_out_and_8_cse & IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse & (~
        (mux_305_nl)) ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0,
          IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0,
          {and_dcpl_236 , and_dcpl_239 , and_dcpl_243});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm <= 1'b0;
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm <= 1'b0;
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_and_9_cse ) begin
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0,
          {and_dcpl_236 , and_dcpl_239 , and_dcpl_243});
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0,
          {and_dcpl_236 , and_dcpl_239 , and_dcpl_243});
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm <= MUX1HOT_s_1_3_2(IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0,
          IsNaN_8U_23U_2_nor_2_mx0w0, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0,
          {and_dcpl_236 , and_dcpl_239 , and_dcpl_243});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_4_nor_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_239 | and_328_rgt) & (~ (mux_314_nl)) ) begin
      IsNaN_8U_23U_4_nor_3_itm_2 <= MUX_s_1_2_2(IsNaN_8U_23U_2_nor_3_mx0w0, alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2,
          and_328_rgt);
    end
  end
  assign FpAlu_8U_23U_mux1h_147_nl = MUX1HOT_s_1_4_2((reg_AluIn_data_sva_4_30_0_1_itm[0]),
      (FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1[0]), AluOut_data_0_0_sva_11, (FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1[0]),
      {FpAlu_8U_23U_nor_dfs_6 , FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_equal_tmp_23
      , FpAlu_8U_23U_equal_tmp_29});
  assign alu_loop_op_mux_209_nl = MUX_s_1_2_2((FpAlu_8U_23U_mux1h_147_nl), AluOut_data_2_0_sva_11,
      alu_loop_op_unequal_tmp_8);
  assign FpAlu_8U_23U_mux1h_151_nl = MUX1HOT_s_1_4_2((reg_AluIn_data_sva_4_62_32_1_itm[0]),
      (FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1[0]), AluOut_data_1_0_sva_12, (FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1[0]),
      {FpAlu_8U_23U_nor_dfs_6 , FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_equal_tmp_23
      , FpAlu_8U_23U_equal_tmp_29});
  assign alu_loop_op_mux_210_nl = MUX_s_1_2_2((FpAlu_8U_23U_mux1h_151_nl), AluOut_data_0_0_sva_11,
      alu_loop_op_unequal_tmp_8);
  assign alu_loop_op_mux_212_nl = MUX_s_1_2_2(FpAlu_8U_23U_o_0_lpi_1_dfm_2, AluOut_data_2_0_lpi_1_dfm_3,
      alu_loop_op_unequal_tmp_8);
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_nl = MUX_v_22_2_2((FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1[22:1]),
      (FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1[22:1]), FpAlu_8U_23U_equal_tmp_29);
  assign FpAlu_8U_23U_not_24_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_and_5_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_FpAlu_8U_23U_mux_nl),
      (FpAlu_8U_23U_not_24_nl));
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl = MUX_v_22_2_2((FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1[22:1]),
      (FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1[22:1]), FpAlu_8U_23U_equal_tmp_29);
  assign FpAlu_8U_23U_not_23_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_and_8_nl = MUX_v_22_2_2(22'b0000000000000000000000, (FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl),
      (FpAlu_8U_23U_not_23_nl));
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl = FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13
      + 8'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl = nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_nl = (~(FpAdd_8U_23U_and_tmp_2 | FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8))
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_6_nl = FpAdd_8U_23U_and_tmp_2 & (~ FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8)
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_28_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8 & FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_9_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_11)
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_mux1h_145_nl = MUX1HOT_v_8_6_2(FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13,
      (alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl), 8'b11111110, else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3,
      (FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1[30:23]), (FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1[30:23]),
      {(FpAdd_8U_23U_and_nl) , (FpAdd_8U_23U_and_6_nl) , (FpAdd_8U_23U_and_28_nl)
      , (FpAdd_8U_23U_and_9_nl) , FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_equal_tmp_29});
  assign FpAlu_8U_23U_not_27_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_and_4_nl = MUX_v_8_2_2(8'b00000000, (FpAlu_8U_23U_mux1h_145_nl),
      (FpAlu_8U_23U_not_27_nl));
  assign nor_406_nl = ~(asn_267 | or_996_tmp);
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13
      + 8'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl = nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl[7:0];
  assign FpAdd_8U_23U_and_29_nl = (~(FpAdd_8U_23U_and_1_tmp_3 | FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8))
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_13_nl = FpAdd_8U_23U_and_1_tmp_3 & (~ FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8)
      & FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_30_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8 & FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAdd_8U_23U_and_15_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_11)
      & FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_mux1h_149_nl = MUX1HOT_v_8_6_2(FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13,
      (alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl), 8'b11111110, else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3,
      (FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1[30:23]), (FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1[30:23]),
      {(FpAdd_8U_23U_and_29_nl) , (FpAdd_8U_23U_and_13_nl) , (FpAdd_8U_23U_and_30_nl)
      , (FpAdd_8U_23U_and_15_nl) , FpAlu_8U_23U_equal_tmp_26 , FpAlu_8U_23U_equal_tmp_29});
  assign FpAlu_8U_23U_not_26_nl = ~ FpAlu_8U_23U_equal_tmp_23;
  assign FpAlu_8U_23U_and_7_nl = MUX_v_8_2_2(8'b00000000, (FpAlu_8U_23U_mux1h_149_nl),
      (FpAlu_8U_23U_not_26_nl));
  assign nor_407_nl = ~(asn_267 | or_997_tmp);
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_9, (~ mux_tmp_2), cfg_alu_algo_rsci_d[0]);
  assign mux_19_nl = MUX_s_1_2_2((mux_18_nl), or_tmp_9, cfg_alu_algo_rsci_d[1]);
  assign mux_20_nl = MUX_s_1_2_2(or_tmp_9, (~ mux_tmp_2), cfg_alu_algo_1_sva_st[0]);
  assign mux_21_nl = MUX_s_1_2_2((mux_20_nl), or_tmp_9, or_28_cse);
  assign mux_22_nl = MUX_s_1_2_2((mux_21_nl), (mux_19_nl), nor_6_cse);
  assign mux_23_nl = MUX_s_1_2_2(or_tmp_9, (mux_22_nl), nor_5_cse);
  assign mux_26_nl = MUX_s_1_2_2(or_tmp_15, (~ mux_tmp_10), cfg_alu_algo_rsci_d[0]);
  assign mux_27_nl = MUX_s_1_2_2((mux_26_nl), or_tmp_15, cfg_alu_algo_rsci_d[1]);
  assign mux_28_nl = MUX_s_1_2_2(or_tmp_15, (~ mux_tmp_10), cfg_alu_algo_1_sva_st[0]);
  assign mux_29_nl = MUX_s_1_2_2((mux_28_nl), or_tmp_15, cfg_alu_algo_1_sva_st[1]);
  assign mux_30_nl = MUX_s_1_2_2((mux_29_nl), (mux_27_nl), nor_6_cse);
  assign mux_31_nl = MUX_s_1_2_2(or_tmp_15, (mux_30_nl), nor_5_cse);
  assign nand_18_nl = ~(cfg_alu_bypass_rsc_triosy_obj_bawt & cfg_alu_src_rsc_triosy_obj_bawt
      & cfg_alu_op_rsc_triosy_obj_bawt & cfg_alu_algo_rsc_triosy_obj_bawt & (~ or_tmp_23));
  assign or_43_nl = cfg_alu_bypass_rsci_d | not_tmp_24;
  assign mux_35_nl = MUX_s_1_2_2((~ alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2),
      (or_43_nl), or_1087_cse);
  assign mux_36_nl = MUX_s_1_2_2((~ alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2),
      (mux_35_nl), and_501_cse);
  assign mux_37_nl = MUX_s_1_2_2((mux_36_nl), (nand_18_nl), io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_38_nl = MUX_s_1_2_2(or_tmp_23, (mux_37_nl), main_stage_v_1);
  assign else_AluOp_data_else_AluOp_data_nor_nl = ~((~(io_read_cfg_alu_bypass_rsc_svs_st_1
      | (~ alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2)))
      | and_dcpl_32);
  assign nor_354_nl = ~((z_out_12[49]) | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign nor_355_nl = ~(alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5 | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign mux_58_nl = MUX_s_1_2_2((nor_355_nl), (nor_354_nl), nor_6_cse);
  assign nor_356_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign mux_59_nl = MUX_s_1_2_2((nor_356_nl), (mux_58_nl), or_1087_cse);
  assign nor_351_nl = ~((z_out_13[49]) | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign nor_352_nl = ~(alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5 | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign mux_60_nl = MUX_s_1_2_2((nor_352_nl), (nor_351_nl), nor_6_cse);
  assign nor_353_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2);
  assign mux_61_nl = MUX_s_1_2_2((nor_353_nl), (mux_60_nl), or_1087_cse);
  assign nor_348_nl = ~((z_out_14[49]) | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign nor_349_nl = ~(alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5 | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign mux_62_nl = MUX_s_1_2_2((nor_349_nl), (nor_348_nl), nor_6_cse);
  assign nor_350_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign mux_63_nl = MUX_s_1_2_2((nor_350_nl), (mux_62_nl), or_1087_cse);
  assign nor_345_nl = ~((z_out_15[49]) | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign nor_346_nl = ~(alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5 | (cfg_alu_algo_1_sva_st_23!=2'b10));
  assign mux_64_nl = MUX_s_1_2_2((nor_346_nl), (nor_345_nl), nor_6_cse);
  assign nor_347_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2);
  assign mux_65_nl = MUX_s_1_2_2((nor_347_nl), (mux_64_nl), or_1087_cse);
  assign nor_344_nl = ~((~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3));
  assign mux_66_nl = MUX_s_1_2_2((~ or_tmp_103), main_stage_v_2, or_1087_cse);
  assign mux_67_nl = MUX_s_1_2_2((mux_66_nl), (nor_344_nl), io_read_cfg_alu_bypass_rsc_svs_st_5);
  assign nor_336_nl = ~(nor_33_cse | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10)
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign nor_337_nl = ~((FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49]) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign mux_69_nl = MUX_s_1_2_2((nor_337_nl), (nor_336_nl), alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2);
  assign and_500_nl = ((~ alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp) | alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1)
      & (mux_69_nl);
  assign nor_338_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10)
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_1_lpi_1_dfm_8
      | IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign mux_70_nl = MUX_s_1_2_2((nor_338_nl), (and_500_nl), nor_6_cse);
  assign nor_334_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (mux_70_nl))));
  assign nor_340_nl = ~((~((~ alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2)
      | (~ alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3)
      | (cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 | IsNaN_8U_23U_land_1_lpi_1_dfm_11
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8)) | alu_loop_op_unequal_tmp_8);
  assign nor_342_nl = ~((~((cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_1_lpi_1_dfm_9
      | IsNaN_8U_23U_land_1_lpi_1_dfm_11 | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23
      | io_read_cfg_alu_bypass_rsc_svs_st_7 | FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8))
      | alu_loop_op_unequal_tmp_8);
  assign mux_73_nl = MUX_s_1_2_2((nor_342_nl), (nor_340_nl), FpAdd_8U_23U_and_tmp_2);
  assign nor_339_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | (mux_73_nl));
  assign mux_74_nl = MUX_s_1_2_2((nor_339_nl), (nor_334_nl), or_1087_cse);
  assign nor_326_nl = ~(nor_37_cse | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10)
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign nor_327_nl = ~((FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49]) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign mux_75_nl = MUX_s_1_2_2((nor_327_nl), (nor_326_nl), alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2);
  assign and_499_nl = ((~ alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp) | alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1)
      & (mux_75_nl);
  assign nor_328_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10)
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_8
      | IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign mux_76_nl = MUX_s_1_2_2((nor_328_nl), (and_499_nl), nor_6_cse);
  assign nor_324_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (mux_76_nl))));
  assign nor_330_nl = ~((~((~ alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2)
      | (~ alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3)
      | (cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 | IsNaN_8U_23U_land_2_lpi_1_dfm_11
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8)) | alu_loop_op_unequal_tmp_8);
  assign nor_332_nl = ~((~((cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_2_lpi_1_dfm_9
      | IsNaN_8U_23U_land_2_lpi_1_dfm_11 | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23
      | io_read_cfg_alu_bypass_rsc_svs_st_7 | FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8))
      | alu_loop_op_unequal_tmp_8);
  assign mux_79_nl = MUX_s_1_2_2((nor_332_nl), (nor_330_nl), FpAdd_8U_23U_and_1_tmp_3);
  assign nor_329_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | (mux_79_nl));
  assign mux_80_nl = MUX_s_1_2_2((nor_329_nl), (nor_324_nl), or_1087_cse);
  assign nor_316_nl = ~(nor_41_cse | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10)
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign nor_317_nl = ~((FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49]) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign mux_81_nl = MUX_s_1_2_2((nor_317_nl), (nor_316_nl), alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2);
  assign and_498_nl = ((~ alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp) | alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1)
      & (mux_81_nl);
  assign nor_318_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10)
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_8
      | IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign mux_82_nl = MUX_s_1_2_2((nor_318_nl), (and_498_nl), nor_6_cse);
  assign nor_314_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (mux_82_nl))));
  assign nor_320_nl = ~((~((~ alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2)
      | (~ alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3)
      | (cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 | IsNaN_8U_23U_land_3_lpi_1_dfm_11
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8)) | alu_loop_op_unequal_tmp_8);
  assign nor_322_nl = ~((~((cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_3_lpi_1_dfm_9
      | IsNaN_8U_23U_land_3_lpi_1_dfm_11 | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23
      | io_read_cfg_alu_bypass_rsc_svs_st_7 | FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8))
      | alu_loop_op_unequal_tmp_8);
  assign mux_85_nl = MUX_s_1_2_2((nor_322_nl), (nor_320_nl), FpAdd_8U_23U_and_2_tmp_3);
  assign nor_319_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | (mux_85_nl));
  assign mux_86_nl = MUX_s_1_2_2((nor_319_nl), (nor_314_nl), or_1087_cse);
  assign nor_310_nl = ~(nor_45_cse | (~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign nor_311_nl = ~((FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49]) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10) |
      io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_lpi_1_dfm_8 | IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign mux_87_nl = MUX_s_1_2_2((nor_311_nl), (nor_310_nl), alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2);
  assign and_497_nl = ((~ alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp) | alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1)
      & (mux_87_nl);
  assign nor_312_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7
      | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22 | IsNaN_8U_23U_1_land_lpi_1_dfm_8
      | IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign mux_88_nl = MUX_s_1_2_2((nor_312_nl), (and_497_nl), nor_6_cse);
  assign or_182_nl = (~ alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2) | (~
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3)
      | (cfg_alu_algo_1_sva_st_25!=2'b10) | IsNaN_8U_23U_1_land_lpi_1_dfm_9 | IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign or_962_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_9 | IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign mux_91_nl = MUX_s_1_2_2((or_962_nl), (or_182_nl), FpAdd_8U_23U_and_3_tmp_3);
  assign nor_313_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | FpAdd_8U_23U_is_inf_lpi_1_dfm_8 | (mux_91_nl));
  assign mux_92_nl = MUX_s_1_2_2((nor_313_nl), (mux_88_nl), or_1087_cse);
  assign nor_307_nl = ~((~ alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign nor_308_nl = ~((~ alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st) | (~
      main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign mux_93_nl = MUX_s_1_2_2((nor_308_nl), (nor_307_nl), nor_6_cse);
  assign nor_309_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (cfg_alu_algo_1_sva_st_25[0]) | (~((cfg_alu_algo_1_sva_st_25[1]) & alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2)));
  assign mux_94_nl = MUX_s_1_2_2((nor_309_nl), (mux_93_nl), or_1087_cse);
  assign nor_304_nl = ~((~ alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign nor_305_nl = ~((~ alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st) | (~
      main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign mux_95_nl = MUX_s_1_2_2((nor_305_nl), (nor_304_nl), nor_6_cse);
  assign nor_306_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (cfg_alu_algo_1_sva_st_25[0]) | (~((cfg_alu_algo_1_sva_st_25[1]) & alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2)));
  assign mux_96_nl = MUX_s_1_2_2((nor_306_nl), (mux_95_nl), or_1087_cse);
  assign nor_301_nl = ~((~ alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign nor_302_nl = ~((~ alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st) | (~
      main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign mux_97_nl = MUX_s_1_2_2((nor_302_nl), (nor_301_nl), nor_6_cse);
  assign nor_303_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (cfg_alu_algo_1_sva_st_25[0]) | (~((cfg_alu_algo_1_sva_st_25[1]) & alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2)));
  assign mux_98_nl = MUX_s_1_2_2((nor_303_nl), (mux_97_nl), or_1087_cse);
  assign nor_298_nl = ~((~ alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp) | (~ main_stage_v_3)
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign nor_299_nl = ~((~ alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st) | (~
      main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6 | (cfg_alu_algo_1_sva_st_24!=2'b10));
  assign mux_99_nl = MUX_s_1_2_2((nor_299_nl), (nor_298_nl), nor_6_cse);
  assign nor_300_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (cfg_alu_algo_1_sva_st_25[0]) | (~((cfg_alu_algo_1_sva_st_25[1]) & alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2)));
  assign mux_100_nl = MUX_s_1_2_2((nor_300_nl), (mux_99_nl), or_1087_cse);
  assign or_1100_nl = FpAlu_8U_23U_equal_tmp_23 | FpAlu_8U_23U_equal_tmp_29 | FpAlu_8U_23U_equal_tmp_26
      | alu_loop_op_unequal_tmp_8 | FpAlu_8U_23U_nor_dfs_6;
  assign or_1106_nl = (~(alu_loop_op_unequal_tmp_8 | (~ FpAlu_8U_23U_nor_dfs_6)))
      | or_dcpl_272 | FpAlu_8U_23U_equal_tmp_23;
  assign mux_383_nl = MUX_s_1_2_2((or_1106_nl), (or_1100_nl), asn_267);
  assign or_280_nl = (~ FpAlu_8U_23U_equal_tmp_32) | (~ FpAlu_8U_23U_equal_tmp_29)
      | alu_loop_op_unequal_tmp_8 | io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_127_nl = MUX_s_1_2_2((or_280_nl), or_tmp_261, or_1087_cse);
  assign nor_274_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | FpAlu_8U_23U_equal_tmp_22 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign nor_275_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_9) | IsNaN_8U_23U_land_3_lpi_1_dfm_11);
  assign mux_128_nl = MUX_s_1_2_2((nor_275_nl), (nor_274_nl), or_1087_cse);
  assign nor_272_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | FpAlu_8U_23U_equal_tmp_22 | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign nor_273_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_9) | IsNaN_8U_23U_land_2_lpi_1_dfm_11);
  assign mux_130_nl = MUX_s_1_2_2((nor_273_nl), (nor_272_nl), or_1087_cse);
  assign nor_270_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | FpAlu_8U_23U_equal_tmp_22 | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign nor_271_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_9) | IsNaN_8U_23U_land_1_lpi_1_dfm_11);
  assign mux_131_nl = MUX_s_1_2_2((nor_271_nl), (nor_270_nl), or_1087_cse);
  assign or_299_nl = (~ FpAlu_8U_23U_equal_tmp_26) | io_read_cfg_alu_bypass_rsc_svs_st_7
      | alu_loop_op_unequal_tmp_8 | io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_132_nl = MUX_s_1_2_2((or_299_nl), or_tmp_280, or_1087_cse);
  assign or_301_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ FpAlu_8U_23U_equal_tmp_26) | io_read_cfg_alu_bypass_rsc_svs_st_7 | alu_loop_op_unequal_tmp_8
      | io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_133_nl = MUX_s_1_2_2((or_301_nl), (mux_132_nl), FpAlu_8U_23U_equal_tmp_25);
  assign or_304_nl = (~ FpAlu_8U_23U_equal_tmp_22) | alu_loop_op_unequal_tmp_7 |
      io_read_cfg_alu_bypass_rsc_svs_7 | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~
      main_stage_v_3);
  assign mux_134_nl = MUX_s_1_2_2(or_tmp_218, (or_304_nl), or_1087_cse);
  assign or_307_nl = nor_269_cse | (~ FpAlu_8U_23U_equal_tmp_22) | alu_loop_op_unequal_tmp_7
      | io_read_cfg_alu_bypass_rsc_svs_7 | io_read_cfg_alu_bypass_rsc_svs_st_6 |
      (~ main_stage_v_3);
  assign mux_135_nl = MUX_s_1_2_2((or_307_nl), (mux_134_nl), FpAlu_8U_23U_equal_tmp_23);
  assign or_312_nl = (~ FpAlu_8U_23U_equal_tmp_35) | (~ FpAlu_8U_23U_equal_tmp_32)
      | (~ FpAlu_8U_23U_equal_tmp_29) | io_read_cfg_alu_bypass_rsc_svs_st_7 | alu_loop_op_unequal_tmp_8
      | io_read_cfg_alu_bypass_rsc_svs_8 | (~ main_stage_v_4);
  assign mux_136_nl = MUX_s_1_2_2((or_312_nl), or_tmp_293, or_1087_cse);
  assign nor_267_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | FpAlu_8U_23U_equal_tmp_22 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8) | IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign nor_268_nl = ~((~ main_stage_v_4) | io_read_cfg_alu_bypass_rsc_svs_8 | alu_loop_op_unequal_tmp_8
      | (~ FpAlu_8U_23U_nor_dfs_6) | FpAlu_8U_23U_equal_tmp_23 | io_read_cfg_alu_bypass_rsc_svs_st_7
      | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_9) | IsNaN_8U_23U_land_lpi_1_dfm_11);
  assign mux_137_nl = MUX_s_1_2_2((nor_268_nl), (nor_267_nl), or_1087_cse);
  assign mux_138_nl = MUX_s_1_2_2(or_tmp_218, or_tmp_280, or_1087_cse);
  assign mux_139_nl = MUX_s_1_2_2(or_tmp_224, or_tmp_103, or_1087_cse);
  assign and_218_nl = (~ nor_tmp_144) & and_dcpl_37;
  assign and_220_nl = (~ nor_tmp_144) & main_stage_v_4 & or_1087_cse & (~ io_read_cfg_alu_bypass_rsc_svs_8);
  assign or_1046_nl = main_stage_v_4 | nor_tmp_144;
  assign or_1048_nl = alu_loop_op_unequal_tmp_8 | FpAlu_8U_23U_equal_tmp_23 | FpAlu_8U_23U_nor_dfs_6
      | FpAlu_8U_23U_equal_tmp_26 | FpAlu_8U_23U_equal_tmp_29 | nor_tmp_144;
  assign mux_nl = MUX_s_1_2_2(nor_tmp_144, (or_1048_nl), main_stage_v_4);
  assign mux_361_nl = MUX_s_1_2_2((mux_nl), (or_1046_nl), io_read_cfg_alu_bypass_rsc_svs_8);
  assign and_729_nl = io_read_cfg_alu_bypass_rsc_svs_8 & main_stage_v_4 & (~ nor_tmp_144);
  assign mux_362_nl = MUX_s_1_2_2((and_729_nl), (mux_361_nl), or_1087_cse);
  assign or_333_nl = alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp | or_tmp_315;
  assign and_496_nl = alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp & (~ or_tmp_315);
  assign mux_145_nl = MUX_s_1_2_2((and_496_nl), (or_333_nl), alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st);
  assign or_334_nl = alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp | or_tmp_315;
  assign and_495_nl = alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp & (~ or_tmp_315);
  assign mux_146_nl = MUX_s_1_2_2((and_495_nl), (or_334_nl), alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st);
  assign or_335_nl = alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp | or_tmp_315;
  assign and_494_nl = alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp & (~ or_tmp_315);
  assign mux_147_nl = MUX_s_1_2_2((and_494_nl), (or_335_nl), alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st);
  assign or_336_nl = alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp | or_tmp_315;
  assign and_493_nl = alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp & (~ or_tmp_315);
  assign mux_148_nl = MUX_s_1_2_2((and_493_nl), (or_336_nl), alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st);
  assign nor_263_nl = ~((cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_4
      | (~ FpAlu_8U_23U_nor_dfs_4) | IsNaN_8U_23U_land_1_lpi_1_dfm_9 | (~ main_stage_v_2)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | io_read_cfg_alu_bypass_rsc_svs_6 |
      alu_loop_op_unequal_tmp_6);
  assign mux_149_nl = MUX_s_1_2_2(nor_264_cse, (nor_263_nl), FpAlu_8U_23U_equal_tmp_21);
  assign nor_265_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (FpAlu_8U_23U_equal_tmp_22
      & ((cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 |
      (~ FpAlu_8U_23U_nor_dfs_5) | IsNaN_8U_23U_land_1_lpi_1_dfm_10)));
  assign mux_150_nl = MUX_s_1_2_2((nor_265_nl), (mux_149_nl), or_1087_cse);
  assign nor_260_nl = ~((cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_4
      | (~ FpAlu_8U_23U_nor_dfs_4) | IsNaN_8U_23U_land_2_lpi_1_dfm_9 | (~ main_stage_v_2)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | io_read_cfg_alu_bypass_rsc_svs_6 |
      alu_loop_op_unequal_tmp_6);
  assign mux_151_nl = MUX_s_1_2_2(nor_264_cse, (nor_260_nl), FpAlu_8U_23U_equal_tmp_21);
  assign nor_262_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (FpAlu_8U_23U_equal_tmp_22
      & ((cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 |
      (~ FpAlu_8U_23U_nor_dfs_5) | IsNaN_8U_23U_land_2_lpi_1_dfm_10)));
  assign mux_152_nl = MUX_s_1_2_2((nor_262_nl), (mux_151_nl), or_1087_cse);
  assign nor_257_nl = ~((cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_3_lpi_1_dfm_st_4
      | (~ FpAlu_8U_23U_nor_dfs_4) | IsNaN_8U_23U_land_3_lpi_1_dfm_9 | (~ main_stage_v_2)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | io_read_cfg_alu_bypass_rsc_svs_6 |
      alu_loop_op_unequal_tmp_6);
  assign mux_153_nl = MUX_s_1_2_2(nor_264_cse, (nor_257_nl), FpAlu_8U_23U_equal_tmp_21);
  assign nor_259_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (FpAlu_8U_23U_equal_tmp_22
      & ((cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 |
      (~ FpAlu_8U_23U_nor_dfs_5) | IsNaN_8U_23U_land_3_lpi_1_dfm_10)));
  assign mux_154_nl = MUX_s_1_2_2((nor_259_nl), (mux_153_nl), or_1087_cse);
  assign nor_254_nl = ~((cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_lpi_1_dfm_st_4
      | (~ FpAlu_8U_23U_nor_dfs_4) | IsNaN_8U_23U_land_lpi_1_dfm_9 | (~ main_stage_v_2)
      | io_read_cfg_alu_bypass_rsc_svs_st_5 | io_read_cfg_alu_bypass_rsc_svs_6 |
      alu_loop_op_unequal_tmp_6);
  assign mux_155_nl = MUX_s_1_2_2(nor_264_cse, (nor_254_nl), FpAlu_8U_23U_equal_tmp_21);
  assign nor_256_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (FpAlu_8U_23U_equal_tmp_22
      & ((cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_lpi_1_dfm_st_5 | (~
      FpAlu_8U_23U_nor_dfs_5) | IsNaN_8U_23U_land_lpi_1_dfm_10)));
  assign mux_156_nl = MUX_s_1_2_2((nor_256_nl), (mux_155_nl), or_1087_cse);
  assign nor_252_nl = ~((z_out_12[49]) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347);
  assign or_961_nl = (~ (z_out_12[49])) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347;
  assign mux_157_nl = MUX_s_1_2_2((or_961_nl), (nor_252_nl), alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm);
  assign nor_251_nl = ~((z_out_13[49]) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347);
  assign or_960_nl = (~ (z_out_13[49])) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347;
  assign mux_158_nl = MUX_s_1_2_2((or_960_nl), (nor_251_nl), alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm);
  assign nor_250_nl = ~((z_out_14[49]) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347);
  assign or_959_nl = (~ (z_out_14[49])) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347;
  assign mux_159_nl = MUX_s_1_2_2((or_959_nl), (nor_250_nl), alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm);
  assign nor_249_nl = ~((z_out_15[49]) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347);
  assign or_958_nl = (~ (z_out_15[49])) | (cfg_alu_algo_1_sva_st_23!=2'b10) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | or_tmp_347;
  assign mux_160_nl = MUX_s_1_2_2((or_958_nl), (nor_249_nl), alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm);
  assign or_400_nl = (cfg_alu_algo_rsci_d!=2'b01);
  assign mux_171_nl = MUX_s_1_2_2((or_400_nl), or_tmp_382, and_489_cse);
  assign mux_172_nl = MUX_s_1_2_2(or_tmp_382, (mux_171_nl), nor_71_cse);
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_nl = (AluOut_data_0_0_sva_9
      & (~ alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1)) | alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign or_422_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | mux_tmp_164;
  assign or_420_nl = (~ FpAlu_8U_23U_equal_tmp_21) | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign mux_181_nl = MUX_s_1_2_2(mux_tmp_165, (or_422_nl), or_420_nl);
  assign mux_182_nl = MUX_s_1_2_2((mux_181_nl), mux_tmp_165, alu_loop_op_unequal_tmp_6);
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_3_nl = (FpAlu_8U_23U_mux1h_33_itm_2
      & (~ alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1)) | alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_2_nl = (FpAlu_8U_23U_mux1h_152_itm_2
      & (~ alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1)) | alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_1_nl = (AluOut_data_1_0_sva_10
      & (~ alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1)) | alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  assign or_438_nl = or_tmp_409 | or_tmp_416;
  assign mux_189_nl = MUX_s_1_2_2((or_438_nl), mux_tmp_173, FpAlu_8U_23U_equal_tmp_25);
  assign or_440_nl = (~ FpAlu_8U_23U_equal_tmp_25) | (~ reg_chn_alu_out_rsci_ld_core_psct_cse)
      | chn_alu_out_rsci_bawt | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7
      | io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ main_stage_v_3);
  assign mux_190_nl = MUX_s_1_2_2((or_440_nl), (mux_189_nl), FpAlu_8U_23U_equal_tmp_24);
  assign or_446_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ FpAlu_8U_23U_equal_tmp_34) | (~ FpAlu_8U_23U_equal_tmp_31) | (~ FpAlu_8U_23U_equal_tmp_28)
      | alu_loop_op_unequal_tmp_7 | io_read_cfg_alu_bypass_rsc_svs_7 | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (~ main_stage_v_3);
  assign mux_193_nl = MUX_s_1_2_2(or_tmp_293, or_tmp_395, or_1087_cse);
  assign or_444_nl = alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_equal_tmp_33) |
      (~ FpAlu_8U_23U_equal_tmp_30) | (~ FpAlu_8U_23U_equal_tmp_27) | io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign mux_194_nl = MUX_s_1_2_2((mux_193_nl), (or_446_nl), or_444_nl);
  assign mux_195_nl = MUX_s_1_2_2(or_tmp_261, or_tmp_395, or_1087_cse);
  assign or_450_nl = (~ reg_chn_alu_out_rsci_ld_core_psct_cse) | chn_alu_out_rsci_bawt
      | (~ FpAlu_8U_23U_equal_tmp_31) | (~ FpAlu_8U_23U_equal_tmp_28) | alu_loop_op_unequal_tmp_7
      | io_read_cfg_alu_bypass_rsc_svs_7 | (~ main_stage_v_3);
  assign nor_80_nl = ~(alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_equal_tmp_30)
      | (~ FpAlu_8U_23U_equal_tmp_27));
  assign mux_196_nl = MUX_s_1_2_2((or_450_nl), (mux_195_nl), nor_80_nl);
  assign nor_237_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ FpAlu_8U_23U_nor_dfs_4)
      | FpAlu_8U_23U_equal_tmp_21 | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7) | IsNaN_8U_23U_land_3_lpi_1_dfm_9
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6);
  assign mux_199_nl = MUX_s_1_2_2((nor_237_nl), nor_236_cse, alu_loop_op_unequal_tmp_6);
  assign nor_238_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | IsNaN_8U_23U_land_3_lpi_1_dfm_10)))));
  assign mux_200_nl = MUX_s_1_2_2((nor_238_nl), (mux_199_nl), or_1087_cse);
  assign nor_232_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ FpAlu_8U_23U_nor_dfs_4)
      | FpAlu_8U_23U_equal_tmp_21 | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7) | IsNaN_8U_23U_land_lpi_1_dfm_9
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6);
  assign mux_203_nl = MUX_s_1_2_2((nor_232_nl), nor_236_cse, alu_loop_op_unequal_tmp_6);
  assign nor_233_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8) | IsNaN_8U_23U_land_lpi_1_dfm_10)))));
  assign mux_204_nl = MUX_s_1_2_2((nor_233_nl), (mux_203_nl), or_1087_cse);
  assign nor_227_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ FpAlu_8U_23U_nor_dfs_4)
      | FpAlu_8U_23U_equal_tmp_21 | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) | IsNaN_8U_23U_land_2_lpi_1_dfm_9
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6);
  assign mux_205_nl = MUX_s_1_2_2((nor_227_nl), nor_236_cse, alu_loop_op_unequal_tmp_6);
  assign nor_228_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | IsNaN_8U_23U_land_2_lpi_1_dfm_10)))));
  assign mux_206_nl = MUX_s_1_2_2((nor_228_nl), (mux_205_nl), or_1087_cse);
  assign nor_222_nl = ~(io_read_cfg_alu_bypass_rsc_svs_st_5 | (~ FpAlu_8U_23U_nor_dfs_4)
      | FpAlu_8U_23U_equal_tmp_21 | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7) | IsNaN_8U_23U_land_1_lpi_1_dfm_9
      | (~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6);
  assign mux_207_nl = MUX_s_1_2_2((nor_222_nl), nor_236_cse, alu_loop_op_unequal_tmp_6);
  assign nor_223_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_7 | (~(alu_loop_op_unequal_tmp_7
      | (~(io_read_cfg_alu_bypass_rsc_svs_st_6 | (~ FpAlu_8U_23U_nor_dfs_5) | FpAlu_8U_23U_equal_tmp_22
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | IsNaN_8U_23U_land_1_lpi_1_dfm_10)))));
  assign mux_208_nl = MUX_s_1_2_2((nor_223_nl), (mux_207_nl), or_1087_cse);
  assign FpAlu_8U_23U_and_9_nl = FpAlu_8U_23U_mux1h_152_itm_2 & (~ FpAlu_8U_23U_equal_tmp_21);
  assign FpAlu_8U_23U_and_nl = FpAlu_8U_23U_mux1h_33_itm_2 & (~ FpAlu_8U_23U_equal_tmp_21);
  assign nor_219_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 |
      io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_nor_dfs_4)
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_7) | IsNaN_8U_23U_land_1_lpi_1_dfm_9);
  assign nor_220_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 |
      io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | (~ IsNaN_8U_23U_1_land_1_lpi_1_dfm_8) | IsNaN_8U_23U_land_1_lpi_1_dfm_10);
  assign mux_209_nl = MUX_s_1_2_2((nor_220_nl), (nor_219_nl), or_1087_cse);
  assign nor_217_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 |
      io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_nor_dfs_4)
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_7) | IsNaN_8U_23U_land_2_lpi_1_dfm_9);
  assign nor_218_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 |
      io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | (~ IsNaN_8U_23U_1_land_2_lpi_1_dfm_8) | IsNaN_8U_23U_land_2_lpi_1_dfm_10);
  assign mux_210_nl = MUX_s_1_2_2((nor_218_nl), (nor_217_nl), or_1087_cse);
  assign nor_215_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 |
      io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_nor_dfs_4)
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_7) | IsNaN_8U_23U_land_3_lpi_1_dfm_9);
  assign nor_216_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 |
      io_read_cfg_alu_bypass_rsc_svs_7 | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5)
      | (~ IsNaN_8U_23U_1_land_3_lpi_1_dfm_8) | IsNaN_8U_23U_land_3_lpi_1_dfm_10);
  assign mux_211_nl = MUX_s_1_2_2((nor_216_nl), (nor_215_nl), or_1087_cse);
  assign nor_213_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | (cfg_alu_algo_1_sva_st_23!=2'b10) | IsNaN_8U_23U_land_lpi_1_dfm_st_4 | io_read_cfg_alu_bypass_rsc_svs_6
      | alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_nor_dfs_4) | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_7)
      | IsNaN_8U_23U_land_lpi_1_dfm_9);
  assign nor_214_nl = ~((~ main_stage_v_3) | io_read_cfg_alu_bypass_rsc_svs_st_6
      | (cfg_alu_algo_1_sva_st_24!=2'b10) | IsNaN_8U_23U_land_lpi_1_dfm_st_5 | io_read_cfg_alu_bypass_rsc_svs_7
      | alu_loop_op_unequal_tmp_7 | (~ FpAlu_8U_23U_nor_dfs_5) | (~ IsNaN_8U_23U_1_land_lpi_1_dfm_8)
      | IsNaN_8U_23U_land_lpi_1_dfm_10);
  assign mux_212_nl = MUX_s_1_2_2((nor_214_nl), (nor_213_nl), or_1087_cse);
  assign FpAlu_8U_23U_or_145_nl = ((~ FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0)
      & FpAlu_8U_23U_and_52_m1c) | (IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 & FpAlu_8U_23U_and_36_m1c);
  assign FpAlu_8U_23U_or_146_nl = (FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0
      & FpAlu_8U_23U_and_52_m1c) | (IsNaN_8U_23U_land_1_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0);
  assign FpAlu_8U_23U_mux1h_144_nl = MUX1HOT_s_1_4_2((else_AluOp_data_0_lpi_1_dfm_mx0[31]),
      (AluIn_data_sva_127[31]), (FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0[31]), (FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0[31]),
      {(FpAlu_8U_23U_or_145_nl) , (FpAlu_8U_23U_or_146_nl) , FpAlu_8U_23U_equal_tmp_mx0w0
      , FpAlu_8U_23U_equal_tmp_2_mx0w0});
  assign FpAlu_8U_23U_or_147_nl = ((~ FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0)
      & FpAlu_8U_23U_and_56_m1c) | (IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 & FpAlu_8U_23U_and_38_m1c);
  assign FpAlu_8U_23U_or_148_nl = (FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0
      & FpAlu_8U_23U_and_56_m1c) | (IsNaN_8U_23U_land_2_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0);
  assign FpAlu_8U_23U_mux1h_148_nl = MUX1HOT_s_1_4_2((else_AluOp_data_1_lpi_1_dfm_mx0[31]),
      (AluIn_data_sva_127[63]), (FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0[31]), (FpCmp_8U_23U_false_o_2_lpi_1_dfm_2[31]),
      {(FpAlu_8U_23U_or_147_nl) , (FpAlu_8U_23U_or_148_nl) , FpAlu_8U_23U_equal_tmp_mx0w0
      , FpAlu_8U_23U_equal_tmp_2_mx0w0});
  assign nor_207_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_equal_tmp_21));
  assign mux_218_nl = MUX_s_1_2_2((nor_207_nl), and_481_cse, or_1087_cse);
  assign nor_206_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6
      | (~ FpAlu_8U_23U_equal_tmp_21));
  assign mux_219_nl = MUX_s_1_2_2((nor_206_nl), and_481_cse, or_1087_cse);
  assign alu_loop_op_else_mux_1_nl = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_1_mx0w0,
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign AluOut_data_or_1_nl = and_dcpl_207 | ((alu_loop_op_else_mux_1_nl) & and_dcpl_208);
  assign alu_loop_op_else_mux_2_nl = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_2_mx0w0,
      IsNaN_8U_23U_4_nor_3_itm_3, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign AluOut_data_or_2_nl = AluOut_data_and_5_cse | ((alu_loop_op_else_mux_2_nl)
      & and_dcpl_208);
  assign alu_loop_op_else_mux_nl = MUX_s_1_2_2(alu_loop_op_else_equal_tmp_2, alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign AluOut_data_and_7_nl = (alu_loop_op_else_mux_nl) & and_dcpl_208;
  assign FpAlu_8U_23U_mux_21_nl = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_1_mx0w0, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign AluOut_data_or_nl = and_dcpl_207 | ((FpAlu_8U_23U_mux_21_nl) & and_dcpl_208);
  assign FpAlu_8U_23U_mux_20_nl = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_2_mx0w0, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign AluOut_data_or_3_nl = AluOut_data_and_5_cse | ((FpAlu_8U_23U_mux_20_nl)
      & and_dcpl_208);
  assign alu_loop_op_else_mux_3_nl = MUX_s_1_2_2(alu_loop_op_else_equal_tmp_2, IsNaN_8U_23U_4_nor_2_itm_2,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign AluOut_data_and_3_nl = (alu_loop_op_else_mux_3_nl) & and_dcpl_208;
  assign nor_203_nl = ~((~ main_stage_v_2) | io_read_cfg_alu_bypass_rsc_svs_st_5
      | io_read_cfg_alu_bypass_rsc_svs_6 | alu_loop_op_unequal_tmp_6 | (~ FpAlu_8U_23U_equal_tmp_24));
  assign mux_223_nl = MUX_s_1_2_2((nor_203_nl), nor_201_cse, or_1087_cse);
  assign nor_195_nl = ~(nor_202_cse | (cfg_precision!=2'b10) | (~ main_stage_v_1)
      | io_read_cfg_alu_bypass_rsc_svs_st_1 | (cfg_alu_algo_1_sva_st_22!=2'b01) |
      (~ cfg_alu_bypass_rsc_triosy_obj_bawt) | (~ cfg_alu_src_rsc_triosy_obj_bawt)
      | (~ cfg_alu_op_rsc_triosy_obj_bawt) | (~ cfg_alu_algo_rsc_triosy_obj_bawt)
      | io_read_cfg_alu_bypass_rsc_svs_5);
  assign mux_225_nl = MUX_s_1_2_2(nor_197_cse, (nor_195_nl), or_1087_cse);
  assign nor_192_nl = ~(nor_202_cse | (cfg_precision!=2'b10) | (~ main_stage_v_1)
      | io_read_cfg_alu_bypass_rsc_svs_st_1 | (cfg_alu_algo_1_sva_st_22!=2'b01) |
      (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01) | (~ cfg_alu_bypass_rsc_triosy_obj_bawt)
      | (~ cfg_alu_src_rsc_triosy_obj_bawt) | (~ cfg_alu_op_rsc_triosy_obj_bawt)
      | (~ cfg_alu_algo_rsc_triosy_obj_bawt) | io_read_cfg_alu_bypass_rsc_svs_5);
  assign mux_226_nl = MUX_s_1_2_2(nor_264_cse, (nor_192_nl), or_1087_cse);
  assign mux_363_nl = MUX_s_1_2_2(or_1055_cse, alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2,
      or_1050_cse);
  assign mux_364_nl = MUX_s_1_2_2(or_1055_cse, alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2,
      or_1050_cse);
  assign or_1069_nl = (cfg_alu_algo_1_sva_2!=2'b01) | (cfg_alu_algo_1_sva_st_22!=2'b01);
  assign mux_365_nl = MUX_s_1_2_2((or_1069_nl), alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2,
      or_1050_cse);
  assign or_1076_nl = (cfg_alu_algo_1_sva_2!=2'b01) | (cfg_alu_algo_1_sva_st_22!=2'b01)
      | (reg_cfg_alu_algo_1_sva_st_13_cse!=2'b01);
  assign mux_366_nl = MUX_s_1_2_2((or_1076_nl), alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2,
      or_1050_cse);
  assign FpAlu_8U_23U_and_74_nl = (((~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0)
      & FpAlu_8U_23U_and_40_m1c) | (IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 & FpAlu_8U_23U_and_24_m1c))
      & and_dcpl_207;
  assign FpAlu_8U_23U_and_75_nl = ((FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0
      & FpAlu_8U_23U_and_40_m1c) | (IsNaN_8U_23U_land_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0))
      & and_dcpl_207;
  assign FpAlu_8U_23U_and_76_nl = FpAlu_8U_23U_equal_tmp_mx0w0 & and_dcpl_207;
  assign FpAlu_8U_23U_and_77_nl = FpAlu_8U_23U_equal_tmp_2_mx0w0 & and_dcpl_207;
  assign alu_loop_op_else_mux_5_nl = MUX_s_1_2_2(FpAlu_8U_23U_equal_tmp_1_mx0w0,
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign FpAlu_8U_23U_and_80_nl = (alu_loop_op_else_mux_5_nl) & and_dcpl_214;
  assign alu_loop_op_else_mux_4_nl = MUX_s_1_2_2(alu_loop_op_else_equal_tmp_2, IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign FpAlu_8U_23U_and_81_nl = (alu_loop_op_else_mux_4_nl) & and_dcpl_214;
  assign FpAlu_8U_23U_and_66_nl = (((~ FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0)
      & FpAlu_8U_23U_and_48_m1c) | (IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 & FpAlu_8U_23U_and_34_m1c))
      & and_297_m1c;
  assign FpAlu_8U_23U_and_67_nl = ((FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0
      & FpAlu_8U_23U_and_48_m1c) | (IsNaN_8U_23U_land_3_lpi_1_dfm_8 & FpAlu_8U_23U_nor_dfs_mx0w0))
      & and_297_m1c;
  assign FpAlu_8U_23U_and_68_nl = FpAlu_8U_23U_equal_tmp_mx0w0 & and_297_m1c;
  assign FpAlu_8U_23U_and_69_nl = FpAlu_8U_23U_equal_tmp_2_mx0w0 & and_297_m1c;
  assign FpAlu_8U_23U_and_72_nl = FpAlu_8U_23U_equal_tmp_1_mx0w0 & and_dcpl_214;
  assign FpAlu_8U_23U_and_73_nl = alu_loop_op_else_equal_tmp_2 & and_dcpl_214;
  assign and_74_nl = or_937_cse & or_tmp_386;
  assign mux_173_nl = MUX_s_1_2_2(nor_tmp_74, (and_74_nl), and_486_cse);
  assign mux_174_nl = MUX_s_1_2_2(or_tmp_386, (mux_173_nl), main_stage_v_1);
  assign nand_30_nl = ~(main_stage_v_1 & (~ nor_tmp_74));
  assign mux_175_nl = MUX_s_1_2_2((nand_30_nl), (mux_174_nl), or_1087_cse);
  assign mux_271_nl = MUX_s_1_2_2(or_tmp_597, or_tmp_596, and_486_cse);
  assign mux_272_nl = MUX_s_1_2_2(or_tmp_597, or_tmp_596, and_501_cse);
  assign or_624_nl = (~((cfg_precision!=2'b10) | cfg_alu_bypass_rsci_d | (~ chn_alu_in_rsci_bawt)))
      | (cfg_alu_algo_1_sva_st[1]) | not_tmp_259;
  assign mux_273_nl = MUX_s_1_2_2(not_tmp_261, (or_624_nl), or_1087_cse);
  assign mux_274_nl = MUX_s_1_2_2(not_tmp_261, (mux_273_nl), and_501_cse);
  assign or_619_nl = (cfg_alu_algo_1_sva_st_22!=2'b01) | (cfg_alu_algo_1_sva_2!=2'b01)
      | io_read_cfg_alu_bypass_rsc_svs_5;
  assign mux_275_nl = MUX_s_1_2_2((mux_274_nl), (mux_272_nl), or_619_nl);
  assign mux_276_nl = MUX_s_1_2_2((mux_275_nl), (mux_271_nl), io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_277_nl = MUX_s_1_2_2(or_tmp_596, (mux_276_nl), main_stage_v_1);
  assign mux_284_nl = MUX_s_1_2_2(mux_tmp_268, mux_tmp_265, and_501_cse);
  assign mux_285_nl = MUX_s_1_2_2((mux_284_nl), mux_281_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_286_nl = MUX_s_1_2_2(mux_tmp_265, (mux_285_nl), main_stage_v_1);
  assign nor_178_nl = ~(and_501_cse | mux_tmp_268);
  assign mux_287_nl = MUX_s_1_2_2((nor_178_nl), nor_177_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nand_35_nl = ~(main_stage_v_1 & (mux_287_nl));
  assign mux_288_nl = MUX_s_1_2_2((nand_35_nl), (mux_286_nl), nor_5_cse);
  assign mux_289_nl = MUX_s_1_2_2(mux_tmp_268, io_read_cfg_alu_bypass_rsc_svs_5,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nand_36_nl = ~(main_stage_v_1 & (~ (mux_289_nl)));
  assign mux_290_nl = MUX_s_1_2_2((nand_36_nl), (mux_288_nl), or_1087_cse);
  assign mux_297_nl = MUX_s_1_2_2(mux_tmp_281, mux_tmp_265, and_501_cse);
  assign mux_298_nl = MUX_s_1_2_2((mux_297_nl), mux_281_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign mux_299_nl = MUX_s_1_2_2(mux_tmp_265, (mux_298_nl), main_stage_v_1);
  assign nor_176_nl = ~(and_501_cse | mux_tmp_281);
  assign mux_300_nl = MUX_s_1_2_2((nor_176_nl), nor_177_cse, io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nand_37_nl = ~(main_stage_v_1 & (mux_300_nl));
  assign mux_301_nl = MUX_s_1_2_2((nand_37_nl), (mux_299_nl), nor_5_cse);
  assign mux_302_nl = MUX_s_1_2_2(mux_tmp_281, io_read_cfg_alu_bypass_rsc_svs_5,
      io_read_cfg_alu_bypass_rsc_svs_st_1);
  assign nand_38_nl = ~(main_stage_v_1 & (~ (mux_302_nl)));
  assign mux_303_nl = MUX_s_1_2_2((nand_38_nl), (mux_301_nl), or_1087_cse);
  assign mux_304_nl = MUX_s_1_2_2(and_451_cse, nor_tmp_126, and_489_cse);
  assign mux_305_nl = MUX_s_1_2_2(nor_tmp_126, (mux_304_nl), nor_71_cse);
  assign mux_313_nl = MUX_s_1_2_2(mux_312_cse, mux_tmp_296, and_489_cse);
  assign mux_314_nl = MUX_s_1_2_2(mux_tmp_296, (mux_313_nl), nor_71_cse);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_15_nl = MUX_v_8_2_2((AluIn_data_sva_127[126:119]),
      (else_AluOp_data_3_lpi_1_dfm_mx0[30:23]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_16_nl = MUX_v_8_2_2((~ (else_AluOp_data_3_lpi_1_dfm_mx0[30:23])),
      (~ (AluIn_data_sva_127[126:119])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp);
  assign nl_acc_4_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_15_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_16_nl)
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[8:0];
  assign z_out_4 = readslicef_9_8_1((acc_4_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_17_nl = MUX_v_8_2_2((AluIn_data_sva_127[94:87]),
      (else_AluOp_data_2_lpi_1_dfm_mx0[30:23]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_18_nl = MUX_v_8_2_2((~ (else_AluOp_data_2_lpi_1_dfm_mx0[30:23])),
      (~ (AluIn_data_sva_127[94:87])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1);
  assign nl_acc_5_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_17_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_18_nl)
      , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[8:0];
  assign z_out_5 = readslicef_9_8_1((acc_5_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_19_nl = MUX_v_8_2_2((AluIn_data_sva_127[62:55]),
      (else_AluOp_data_1_lpi_1_dfm_mx2_30_0[30:23]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_20_nl = MUX_v_8_2_2((~ (else_AluOp_data_1_lpi_1_dfm_mx2_30_0[30:23])),
      (~ (AluIn_data_sva_127[62:55])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2);
  assign nl_acc_6_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_19_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_20_nl)
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[8:0];
  assign z_out_6 = readslicef_9_8_1((acc_6_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_21_nl = MUX_v_8_2_2((AluIn_data_sva_127[30:23]),
      (else_AluOp_data_0_lpi_1_dfm_mx0[30:23]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_22_nl = MUX_v_8_2_2((~ (else_AluOp_data_0_lpi_1_dfm_mx0[30:23])),
      (~ (AluIn_data_sva_127[30:23])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3);
  assign nl_acc_7_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_21_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_22_nl)
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[8:0];
  assign z_out_7 = readslicef_9_8_1((acc_7_nl));
  assign FpAdd_8U_23U_else_2_mux_8_nl = MUX_v_49_2_2((~ FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0),
      FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp);
  assign FpAdd_8U_23U_else_2_mux_9_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0,
      FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp);
  assign nl_acc_12_nl = ({(~ FpAdd_8U_23U_if_2_and_tmp) , (FpAdd_8U_23U_else_2_mux_8_nl)
      , (~ FpAdd_8U_23U_if_2_and_tmp)}) + conv_u2u_50_51({(FpAdd_8U_23U_else_2_mux_9_nl)
      , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[50:0];
  assign z_out_12 = readslicef_51_50_1((acc_12_nl));
  assign FpAdd_8U_23U_else_2_mux_10_nl = MUX_v_49_2_2((~ FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0),
      FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp_1);
  assign FpAdd_8U_23U_else_2_mux_11_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0,
      FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp_1);
  assign nl_acc_13_nl = ({(~ FpAdd_8U_23U_if_2_and_tmp_1) , (FpAdd_8U_23U_else_2_mux_10_nl)
      , (~ FpAdd_8U_23U_if_2_and_tmp_1)}) + conv_u2u_50_51({(FpAdd_8U_23U_else_2_mux_11_nl)
      , 1'b1});
  assign acc_13_nl = nl_acc_13_nl[50:0];
  assign z_out_13 = readslicef_51_50_1((acc_13_nl));
  assign FpAdd_8U_23U_else_2_mux_12_nl = MUX_v_49_2_2((~ FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0),
      FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp_2);
  assign FpAdd_8U_23U_else_2_mux_13_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0,
      FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp_2);
  assign nl_acc_14_nl = ({(~ FpAdd_8U_23U_if_2_and_tmp_2) , (FpAdd_8U_23U_else_2_mux_12_nl)
      , (~ FpAdd_8U_23U_if_2_and_tmp_2)}) + conv_u2u_50_51({(FpAdd_8U_23U_else_2_mux_13_nl)
      , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[50:0];
  assign z_out_14 = readslicef_51_50_1((acc_14_nl));
  assign FpAdd_8U_23U_else_2_mux_14_nl = MUX_v_49_2_2((~ FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0),
      FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp_3);
  assign FpAdd_8U_23U_else_2_mux_15_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0,
      FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0, FpAdd_8U_23U_if_2_and_tmp_3);
  assign nl_acc_15_nl = ({(~ FpAdd_8U_23U_if_2_and_tmp_3) , (FpAdd_8U_23U_else_2_mux_14_nl)
      , (~ FpAdd_8U_23U_if_2_and_tmp_3)}) + conv_u2u_50_51({(FpAdd_8U_23U_else_2_mux_15_nl)
      , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[50:0];
  assign z_out_15 = readslicef_51_50_1((acc_15_nl));

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function [21:0] MUX1HOT_v_22_3_2;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [2:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    MUX1HOT_v_22_3_2 = result;
  end
  endfunction


  function [21:0] MUX1HOT_v_22_4_2;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [3:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    MUX1HOT_v_22_4_2 = result;
  end
  endfunction


  function [30:0] MUX1HOT_v_31_3_2;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [2:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | ( input_1 & {31{sel[1]}});
    result = result | ( input_2 & {31{sel[2]}});
    MUX1HOT_v_31_3_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_7_2;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [6:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    MUX1HOT_v_8_7_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [48:0] MUX_v_49_2_2;
    input [48:0] input_0;
    input [48:0] input_1;
    input [0:0] sel;
    reg [48:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_49_2_2 = result;
  end
  endfunction


  function [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_24_1_23;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 23;
    readslicef_24_1_23 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function [49:0] readslicef_51_50_1;
    input [50:0] vector;
    reg [50:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_51_50_1 = tmp[49:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function [31:0] signext_32_31;
    input [30:0] vector;
  begin
    signext_32_31= {{1{vector[30]}}, vector};
  end
  endfunction


  function  [32:0] conv_s2s_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2s_32_33 = {vector[31], vector};
  end
  endfunction


  function  [2:0] conv_s2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction


  function  [8:0] conv_s2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_9 = {vector[7], vector};
  end
  endfunction


  function  [33:0] conv_s2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_s2u_33_34 = {vector[32], vector};
  end
  endfunction


  function  [8:0] conv_u2s_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function  [22:0] conv_u2u_1_23 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction


  function  [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function  [23:0] conv_u2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_u2u_23_24 = {1'b0, vector};
  end
  endfunction


  function  [50:0] conv_u2u_50_51 ;
    input [49:0]  vector ;
  begin
    conv_u2u_50_51 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_mul
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_mul (
  nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_z, chn_mul_in_rsc_vz, chn_mul_in_rsc_lz,
      chn_mul_op_rsc_z, chn_mul_op_rsc_vz, chn_mul_op_rsc_lz, cfg_mul_bypass_rsc_z,
      cfg_mul_bypass_rsc_triosy_lz, cfg_mul_prelu_rsc_z, cfg_mul_prelu_rsc_triosy_lz,
      cfg_mul_src_rsc_z, cfg_mul_src_rsc_triosy_lz, cfg_mul_op_rsc_z, cfg_mul_op_rsc_triosy_lz,
      cfg_truncate_rsc_z, cfg_truncate_rsc_triosy_lz, cfg_precision, chn_mul_out_rsc_z,
      chn_mul_out_rsc_vz, chn_mul_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_mul_in_rsc_z;
  input chn_mul_in_rsc_vz;
  output chn_mul_in_rsc_lz;
  input [127:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  input cfg_mul_bypass_rsc_z;
  output cfg_mul_bypass_rsc_triosy_lz;
  input cfg_mul_prelu_rsc_z;
  output cfg_mul_prelu_rsc_triosy_lz;
  input cfg_mul_src_rsc_z;
  output cfg_mul_src_rsc_triosy_lz;
  input [31:0] cfg_mul_op_rsc_z;
  output cfg_mul_op_rsc_triosy_lz;
  input [9:0] cfg_truncate_rsc_z;
  output cfg_truncate_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [127:0] chn_mul_out_rsc_z;
  input chn_mul_out_rsc_vz;
  output chn_mul_out_rsc_lz;


  // Interconnect Declarations
  wire chn_mul_in_rsci_oswt;
  wire chn_mul_in_rsci_oswt_unreg;
  wire chn_mul_op_rsci_oswt;
  wire chn_mul_op_rsci_oswt_unreg;
  wire cfg_mul_bypass_rsci_d;
  wire cfg_mul_prelu_rsci_d;
  wire cfg_mul_src_rsci_d;
  wire [31:0] cfg_mul_op_rsci_d;
  wire [9:0] cfg_truncate_rsci_d;
  wire chn_mul_out_rsci_oswt;
  wire chn_mul_out_rsci_oswt_unreg;
  wire cfg_mul_bypass_rsc_triosy_obj_oswt;
  wire cfg_mul_prelu_rsc_triosy_obj_oswt;
  wire cfg_mul_src_rsc_triosy_obj_oswt;
  wire cfg_mul_op_rsc_triosy_obj_oswt;
  wire cfg_truncate_rsc_triosy_obj_oswt;
  wire cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd1)) cfg_mul_bypass_rsci (
      .d(cfg_mul_bypass_rsci_d),
      .z(cfg_mul_bypass_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd4),
  .width(32'sd1)) cfg_mul_prelu_rsci (
      .d(cfg_mul_prelu_rsci_d),
      .z(cfg_mul_prelu_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd5),
  .width(32'sd1)) cfg_mul_src_rsci (
      .d(cfg_mul_src_rsci_d),
      .z(cfg_mul_src_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd6),
  .width(32'sd32)) cfg_mul_op_rsci (
      .d(cfg_mul_op_rsci_d),
      .z(cfg_mul_op_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd7),
  .width(32'sd10)) cfg_truncate_rsci (
      .d(cfg_truncate_rsci_d),
      .z(cfg_truncate_rsc_z)
    );
  SDP_Y_CORE_chn_mul_in_rsci_unreg chn_mul_in_rsci_unreg_inst (
      .in_0(chn_mul_in_rsci_oswt_unreg),
      .outsig(chn_mul_in_rsci_oswt)
    );
  SDP_Y_CORE_chn_mul_op_rsci_unreg chn_mul_op_rsci_unreg_inst (
      .in_0(chn_mul_op_rsci_oswt_unreg),
      .outsig(chn_mul_op_rsci_oswt)
    );
  SDP_Y_CORE_chn_mul_out_rsci_unreg chn_mul_out_rsci_unreg_inst (
      .in_0(chn_mul_out_rsci_oswt_unreg),
      .outsig(chn_mul_out_rsci_oswt)
    );
  SDP_Y_CORE_cfg_mul_bypass_rsc_triosy_obj_unreg cfg_mul_bypass_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_bypass_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_mul_prelu_rsc_triosy_obj_unreg cfg_mul_prelu_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_prelu_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_mul_src_rsc_triosy_obj_unreg cfg_mul_src_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_src_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_mul_op_rsc_triosy_obj_unreg cfg_mul_op_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_mul_op_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_truncate_rsc_triosy_obj_unreg cfg_truncate_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_truncate_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_Y_mul_core Y_mul_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsc_z(chn_mul_in_rsc_z),
      .chn_mul_in_rsc_vz(chn_mul_in_rsc_vz),
      .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz),
      .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
      .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
      .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz),
      .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz),
      .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz),
      .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz),
      .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz),
      .cfg_truncate_rsc_triosy_lz(cfg_truncate_rsc_triosy_lz),
      .cfg_precision(cfg_precision),
      .chn_mul_out_rsc_z(chn_mul_out_rsc_z),
      .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz),
      .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz),
      .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
      .chn_mul_in_rsci_oswt_unreg(chn_mul_in_rsci_oswt_unreg),
      .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
      .chn_mul_op_rsci_oswt_unreg(chn_mul_op_rsci_oswt_unreg),
      .cfg_mul_bypass_rsci_d(cfg_mul_bypass_rsci_d),
      .cfg_mul_prelu_rsci_d(cfg_mul_prelu_rsci_d),
      .cfg_mul_src_rsci_d(cfg_mul_src_rsci_d),
      .cfg_mul_op_rsci_d(cfg_mul_op_rsci_d),
      .cfg_truncate_rsci_d(cfg_truncate_rsci_d),
      .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
      .chn_mul_out_rsci_oswt_unreg(chn_mul_out_rsci_oswt_unreg),
      .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
      .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
      .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
      .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
      .cfg_truncate_rsc_triosy_obj_oswt(cfg_truncate_rsc_triosy_obj_oswt),
      .cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff(cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SDP_Y_CORE_Y_alu
// ------------------------------------------------------------------


module SDP_Y_CORE_Y_alu (
  nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz,
      chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, cfg_alu_bypass_rsc_z,
      cfg_alu_bypass_rsc_triosy_lz, cfg_alu_src_rsc_z, cfg_alu_src_rsc_triosy_lz,
      cfg_alu_op_rsc_z, cfg_alu_op_rsc_triosy_lz, cfg_alu_algo_rsc_z, cfg_alu_algo_rsc_triosy_lz,
      cfg_precision, chn_alu_out_rsc_z, chn_alu_out_rsc_vz, chn_alu_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_alu_in_rsc_z;
  input chn_alu_in_rsc_vz;
  output chn_alu_in_rsc_lz;
  input [127:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  input cfg_alu_bypass_rsc_z;
  output cfg_alu_bypass_rsc_triosy_lz;
  input cfg_alu_src_rsc_z;
  output cfg_alu_src_rsc_triosy_lz;
  input [31:0] cfg_alu_op_rsc_z;
  output cfg_alu_op_rsc_triosy_lz;
  input [1:0] cfg_alu_algo_rsc_z;
  output cfg_alu_algo_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [127:0] chn_alu_out_rsc_z;
  input chn_alu_out_rsc_vz;
  output chn_alu_out_rsc_lz;


  // Interconnect Declarations
  wire chn_alu_in_rsci_oswt;
  wire chn_alu_in_rsci_oswt_unreg;
  wire chn_alu_op_rsci_oswt;
  wire chn_alu_op_rsci_oswt_unreg;
  wire cfg_alu_bypass_rsci_d;
  wire cfg_alu_src_rsci_d;
  wire [31:0] cfg_alu_op_rsci_d;
  wire [1:0] cfg_alu_algo_rsci_d;
  wire chn_alu_out_rsci_oswt;
  wire chn_alu_out_rsci_oswt_unreg;
  wire cfg_alu_bypass_rsc_triosy_obj_oswt;
  wire cfg_alu_src_rsc_triosy_obj_oswt;
  wire cfg_alu_op_rsc_triosy_obj_oswt;
  wire cfg_alu_algo_rsc_triosy_obj_oswt;
  wire cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_iff;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd15),
  .width(32'sd1)) cfg_alu_bypass_rsci (
      .d(cfg_alu_bypass_rsci_d),
      .z(cfg_alu_bypass_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd16),
  .width(32'sd1)) cfg_alu_src_rsci (
      .d(cfg_alu_src_rsci_d),
      .z(cfg_alu_src_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd17),
  .width(32'sd32)) cfg_alu_op_rsci (
      .d(cfg_alu_op_rsci_d),
      .z(cfg_alu_op_rsc_z)
    );
  SDP_Y_CORE_mgc_in_wire_v1 #(.rscid(32'sd18),
  .width(32'sd2)) cfg_alu_algo_rsci (
      .d(cfg_alu_algo_rsci_d),
      .z(cfg_alu_algo_rsc_z)
    );
  SDP_Y_CORE_chn_alu_in_rsci_unreg chn_alu_in_rsci_unreg_inst (
      .in_0(chn_alu_in_rsci_oswt_unreg),
      .outsig(chn_alu_in_rsci_oswt)
    );
  SDP_Y_CORE_chn_alu_op_rsci_unreg chn_alu_op_rsci_unreg_inst (
      .in_0(chn_alu_op_rsci_oswt_unreg),
      .outsig(chn_alu_op_rsci_oswt)
    );
  SDP_Y_CORE_chn_alu_out_rsci_unreg chn_alu_out_rsci_unreg_inst (
      .in_0(chn_alu_out_rsci_oswt_unreg),
      .outsig(chn_alu_out_rsci_oswt)
    );
  SDP_Y_CORE_cfg_alu_bypass_rsc_triosy_obj_unreg cfg_alu_bypass_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_bypass_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_alu_src_rsc_triosy_obj_unreg cfg_alu_src_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_src_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_alu_op_rsc_triosy_obj_unreg cfg_alu_op_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_op_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_cfg_alu_algo_rsc_triosy_obj_unreg cfg_alu_algo_rsc_triosy_obj_unreg_inst (
      .in_0(cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_iff),
      .outsig(cfg_alu_algo_rsc_triosy_obj_oswt)
    );
  SDP_Y_CORE_Y_alu_core Y_alu_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsc_z(chn_alu_in_rsc_z),
      .chn_alu_in_rsc_vz(chn_alu_in_rsc_vz),
      .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz),
      .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
      .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
      .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz),
      .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz),
      .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz),
      .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz),
      .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz),
      .cfg_precision(cfg_precision),
      .chn_alu_out_rsc_z(chn_alu_out_rsc_z),
      .chn_alu_out_rsc_vz(chn_alu_out_rsc_vz),
      .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz),
      .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
      .chn_alu_in_rsci_oswt_unreg(chn_alu_in_rsci_oswt_unreg),
      .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
      .chn_alu_op_rsci_oswt_unreg(chn_alu_op_rsci_oswt_unreg),
      .cfg_alu_bypass_rsci_d(cfg_alu_bypass_rsci_d),
      .cfg_alu_src_rsci_d(cfg_alu_src_rsci_d),
      .cfg_alu_op_rsci_d(cfg_alu_op_rsci_d),
      .cfg_alu_algo_rsci_d(cfg_alu_algo_rsci_d),
      .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
      .chn_alu_out_rsci_oswt_unreg(chn_alu_out_rsci_oswt_unreg),
      .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
      .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
      .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
      .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
      .cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff(cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_SDP_CORE_Y_core
// ------------------------------------------------------------------


module NV_NVDLA_SDP_CORE_Y_core (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsc_z, chn_data_in_rsc_vz, chn_data_in_rsc_lz,
      chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, chn_mul_op_rsc_z, chn_mul_op_rsc_vz,
      chn_mul_op_rsc_lz, cfg_alu_bypass_rsc_z, cfg_alu_bypass_rsc_triosy_lz, cfg_alu_src_rsc_z,
      cfg_alu_src_rsc_triosy_lz, cfg_alu_op_rsc_z, cfg_alu_op_rsc_triosy_lz, cfg_alu_algo_rsc_z,
      cfg_alu_algo_rsc_triosy_lz, cfg_mul_bypass_rsc_z, cfg_mul_bypass_rsc_triosy_lz,
      cfg_mul_src_rsc_z, cfg_mul_src_rsc_triosy_lz, cfg_mul_op_rsc_z, cfg_mul_op_rsc_triosy_lz,
      cfg_truncate_rsc_z, cfg_truncate_rsc_triosy_lz, cfg_mul_prelu_rsc_z, cfg_mul_prelu_rsc_triosy_lz,
      cfg_precision, chn_data_out_rsc_z, chn_data_out_rsc_vz, chn_data_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [127:0] chn_data_in_rsc_z;
  input chn_data_in_rsc_vz;
  output chn_data_in_rsc_lz;
  input [127:0] chn_alu_op_rsc_z;
  input chn_alu_op_rsc_vz;
  output chn_alu_op_rsc_lz;
  input [127:0] chn_mul_op_rsc_z;
  input chn_mul_op_rsc_vz;
  output chn_mul_op_rsc_lz;
  input cfg_alu_bypass_rsc_z;
  output cfg_alu_bypass_rsc_triosy_lz;
  input cfg_alu_src_rsc_z;
  output cfg_alu_src_rsc_triosy_lz;
  input [31:0] cfg_alu_op_rsc_z;
  output cfg_alu_op_rsc_triosy_lz;
  input [1:0] cfg_alu_algo_rsc_z;
  output cfg_alu_algo_rsc_triosy_lz;
  input cfg_mul_bypass_rsc_z;
  output cfg_mul_bypass_rsc_triosy_lz;
  input cfg_mul_src_rsc_z;
  output cfg_mul_src_rsc_triosy_lz;
  input [31:0] cfg_mul_op_rsc_z;
  output cfg_mul_op_rsc_triosy_lz;
  input [9:0] cfg_truncate_rsc_z;
  output cfg_truncate_rsc_triosy_lz;
  input cfg_mul_prelu_rsc_z;
  output cfg_mul_prelu_rsc_triosy_lz;
  input [1:0] cfg_precision;
  output [127:0] chn_data_out_rsc_z;
  input chn_data_out_rsc_vz;
  output chn_data_out_rsc_lz;


  // Interconnect Declarations
  wire [127:0] chn_mul_out_rsc_z_nY_mul_inst;
  wire chn_mul_out_rsc_vz_nY_mul_inst;
  wire [127:0] chn_alu_in_rsc_z_nY_alu_inst;
  wire chn_alu_in_rsc_vz_nY_alu_inst;
  wire [127:0] chn_alu_out_rsc_z_nY_alu_inst;
  wire chn_mul_in_rsc_lz_nY_mul_inst_bud;
  wire chn_mul_op_rsc_lz_nY_mul_inst_bud;
  wire cfg_mul_bypass_rsc_triosy_lz_nY_mul_inst_bud;
  wire cfg_mul_prelu_rsc_triosy_lz_nY_mul_inst_bud;
  wire cfg_mul_src_rsc_triosy_lz_nY_mul_inst_bud;
  wire cfg_mul_op_rsc_triosy_lz_nY_mul_inst_bud;
  wire cfg_truncate_rsc_triosy_lz_nY_mul_inst_bud;
  wire chn_mul_out_rsc_lz_nY_mul_inst_bud;
  wire chn_alu_in_rsc_lz_nY_alu_inst_bud;
  wire chn_alu_op_rsc_lz_nY_alu_inst_bud;
  wire cfg_alu_bypass_rsc_triosy_lz_nY_alu_inst_bud;
  wire cfg_alu_src_rsc_triosy_lz_nY_alu_inst_bud;
  wire cfg_alu_op_rsc_triosy_lz_nY_alu_inst_bud;
  wire cfg_alu_algo_rsc_triosy_lz_nY_alu_inst_bud;
  wire chn_alu_out_rsc_lz_nY_alu_inst_bud;
  wire chn_mul_out_unc_2;


  // Interconnect Declarations for Component Instantiations 
  SDP_Y_CORE_mgc_pipe_v10 #(.rscid(32'sd38),
  .width(32'sd128),
  .sz_width(32'sd1),
  .fifo_sz(32'sd5),
  .log2_sz(32'sd3),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) chn_mul_out_cns_pipe (
      .clk(nvdla_core_clk),
      .en(1'b0),
      .arst(nvdla_core_rstn),
      .srst(1'b1),
      .ldin(chn_alu_in_rsc_lz_nY_alu_inst_bud),
      .vdin(chn_alu_in_rsc_vz_nY_alu_inst),
      .din(chn_alu_in_rsc_z_nY_alu_inst),
      .ldout(chn_mul_out_rsc_lz_nY_mul_inst_bud),
      .vdout(chn_mul_out_rsc_vz_nY_mul_inst),
      .dout(chn_mul_out_rsc_z_nY_mul_inst),
      .sd(chn_mul_out_unc_2)
    );
  SDP_Y_CORE_Y_mul Y_mul_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_mul_in_rsc_z(chn_data_in_rsc_z),
      .chn_mul_in_rsc_vz(chn_data_in_rsc_vz),
      .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz_nY_mul_inst_bud),
      .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
      .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
      .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz_nY_mul_inst_bud),
      .cfg_mul_bypass_rsc_z(cfg_mul_bypass_rsc_z),
      .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz_nY_mul_inst_bud),
      .cfg_mul_prelu_rsc_z(cfg_mul_prelu_rsc_z),
      .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz_nY_mul_inst_bud),
      .cfg_mul_src_rsc_z(cfg_mul_src_rsc_z),
      .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz_nY_mul_inst_bud),
      .cfg_mul_op_rsc_z(cfg_mul_op_rsc_z),
      .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz_nY_mul_inst_bud),
      .cfg_truncate_rsc_z(cfg_truncate_rsc_z),
      .cfg_truncate_rsc_triosy_lz(cfg_truncate_rsc_triosy_lz_nY_mul_inst_bud),
      .cfg_precision(cfg_precision),
      .chn_mul_out_rsc_z(chn_mul_out_rsc_z_nY_mul_inst),
      .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz_nY_mul_inst),
      .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz_nY_mul_inst_bud)
    );
  SDP_Y_CORE_Y_alu Y_alu_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_alu_in_rsc_z(chn_alu_in_rsc_z_nY_alu_inst),
      .chn_alu_in_rsc_vz(chn_alu_in_rsc_vz_nY_alu_inst),
      .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz_nY_alu_inst_bud),
      .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
      .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
      .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz_nY_alu_inst_bud),
      .cfg_alu_bypass_rsc_z(cfg_alu_bypass_rsc_z),
      .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz_nY_alu_inst_bud),
      .cfg_alu_src_rsc_z(cfg_alu_src_rsc_z),
      .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz_nY_alu_inst_bud),
      .cfg_alu_op_rsc_z(cfg_alu_op_rsc_z),
      .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz_nY_alu_inst_bud),
      .cfg_alu_algo_rsc_z(cfg_alu_algo_rsc_z),
      .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz_nY_alu_inst_bud),
      .cfg_precision(cfg_precision),
      .chn_alu_out_rsc_z(chn_alu_out_rsc_z_nY_alu_inst),
      .chn_alu_out_rsc_vz(chn_data_out_rsc_vz),
      .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz_nY_alu_inst_bud)
    );
  assign chn_data_in_rsc_lz = chn_mul_in_rsc_lz_nY_mul_inst_bud;
  assign chn_mul_op_rsc_lz = chn_mul_op_rsc_lz_nY_mul_inst_bud;
  assign cfg_mul_bypass_rsc_triosy_lz = cfg_mul_bypass_rsc_triosy_lz_nY_mul_inst_bud;
  assign cfg_mul_prelu_rsc_triosy_lz = cfg_mul_prelu_rsc_triosy_lz_nY_mul_inst_bud;
  assign cfg_mul_src_rsc_triosy_lz = cfg_mul_src_rsc_triosy_lz_nY_mul_inst_bud;
  assign cfg_mul_op_rsc_triosy_lz = cfg_mul_op_rsc_triosy_lz_nY_mul_inst_bud;
  assign cfg_truncate_rsc_triosy_lz = cfg_truncate_rsc_triosy_lz_nY_mul_inst_bud;
  assign chn_alu_op_rsc_lz = chn_alu_op_rsc_lz_nY_alu_inst_bud;
  assign cfg_alu_bypass_rsc_triosy_lz = cfg_alu_bypass_rsc_triosy_lz_nY_alu_inst_bud;
  assign cfg_alu_src_rsc_triosy_lz = cfg_alu_src_rsc_triosy_lz_nY_alu_inst_bud;
  assign cfg_alu_op_rsc_triosy_lz = cfg_alu_op_rsc_triosy_lz_nY_alu_inst_bud;
  assign cfg_alu_algo_rsc_triosy_lz = cfg_alu_algo_rsc_triosy_lz_nY_alu_inst_bud;
  assign chn_data_out_rsc_lz = chn_alu_out_rsc_lz_nY_alu_inst_bud;
  assign chn_data_out_rsc_z = chn_alu_out_rsc_z_nY_alu_inst;
endmodule



